
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RV32I is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RV32I;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RV32I.all;

entity RV32I is

   port( Clk, Rst : in std_logic;  IRAM_DOUT, RF_RD1_DATA, RF_RD2_DATA, 
         DRAM_DOUT : in std_logic_vector (31 downto 0);  IRAM_ADD : out 
         std_logic_vector (31 downto 0);  RF_RD1_EN, RF_RD2_EN, RF_WR_EN : out 
         std_logic;  RF_RD1_ADD, RF_RD2_ADD, RF_WR_ADD : out std_logic_vector 
         (4 downto 0);  RF_WR_DATA : out std_logic_vector (31 downto 0);  
         DRAM_WE, DRAM_RE : out std_logic;  DRAM_ADD, DRAM_DIN : out 
         std_logic_vector (31 downto 0));

end RV32I;

architecture SYN_RV32I_rtl of RV32I is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, RF_RD1_ADD_4_port, 
      RF_RD1_ADD_3_port, RF_RD1_ADD_2_port, RF_RD1_ADD_1_port, 
      RF_RD1_ADD_0_port, RF_RD2_ADD_4_port, RF_RD2_ADD_3_port, 
      RF_RD2_ADD_2_port, RF_RD2_ADD_1_port, RF_RD2_ADD_0_port, DRAM_ADD_31_port
      , DRAM_ADD_30_port, DRAM_ADD_29_port, DRAM_ADD_28_port, DRAM_ADD_27_port,
      DRAM_ADD_26_port, DRAM_ADD_25_port, DRAM_ADD_24_port, DRAM_ADD_23_port, 
      DRAM_ADD_22_port, DRAM_ADD_21_port, DRAM_ADD_20_port, DRAM_ADD_19_port, 
      DRAM_ADD_18_port, DRAM_ADD_17_port, DRAM_ADD_16_port, DRAM_ADD_15_port, 
      DRAM_ADD_14_port, DRAM_ADD_13_port, DRAM_ADD_12_port, DRAM_ADD_11_port, 
      DRAM_ADD_10_port, DRAM_ADD_9_port, DRAM_ADD_8_port, DRAM_ADD_7_port, 
      DRAM_ADD_6_port, DRAM_ADD_5_port, DRAM_ADD_4_port, DRAM_ADD_3_port, 
      DRAM_ADD_2_port, DRAM_ADD_1_port, DRAM_ADD_0_port, PC_SEL_i, IMM_SEL_i, 
      RF_WE_MEM_i, WB_MUX_SEL_MEM_i, BRANCH_EN_i, CU_IxN52, CU_IxN51, 
      CU_Ixcw2_i_10_port, CU_Ixcw2_i_11_port, CU_Ixcw2_i_12_port, 
      CU_Ixcw3_0_port, CU_Ixcw3_1_port, CU_Ixcw3_2_port, CU_Ixcw3_3_port, 
      CU_Ixcw2_0_port, CU_Ixcw2_1_port, CU_Ixcw2_2_port, CU_Ixcw2_3_port, 
      CU_Ixcw2_4_port, CU_Ixcw2_5_port, CU_Ixcw2_6_port, CU_Ixcw1_0_port, 
      CU_Ixcw1_1_port, CU_Ixcw1_2_port, CU_Ixcw1_4_port, CU_Ixcw1_5_port, 
      CU_Ixcw1_6_port, CU_Ixcw1_7_port, CU_Ixcw1_8_port, CU_Ixcw1_9_port, 
      CU_Ixcw1_10_port, CU_Ixcw1_14_port, CU_Ixcw_LUT_0_port, 
      CU_Ixcw_LUT_1_port, CU_Ixcw_LUT_2_port, CU_Ixcw_LUT_4_port, 
      CU_Ixcw_LUT_5_port, CU_Ixcw_LUT_6_port, CU_Ixcw_LUT_7_port, 
      CU_Ixcw_LUT_8_port, CU_Ixcw_LUT_9_port, CU_Ixcw_LUT_10_port, 
      CU_Ixcw_LUT_15_port, CU_Ixcw_LUT_16_port, CU_IxN25, CU_IxN24, CU_IxN23, 
      DATAPATH_IxALUOUT_Data1_0_port, DATAPATH_IxALUOUT_Data1_1_port, 
      DATAPATH_IxALUOUT_Data1_2_port, DATAPATH_IxALUOUT_Data1_3_port, 
      DATAPATH_IxALUOUT_Data1_4_port, DATAPATH_IxALUOUT_Data1_5_port, 
      DATAPATH_IxALUOUT_Data1_6_port, DATAPATH_IxALUOUT_Data1_7_port, 
      DATAPATH_IxALUOUT_Data1_8_port, DATAPATH_IxALUOUT_Data1_9_port, 
      DATAPATH_IxALUOUT_Data1_10_port, DATAPATH_IxALUOUT_Data1_11_port, 
      DATAPATH_IxALUOUT_Data1_12_port, DATAPATH_IxALUOUT_Data1_13_port, 
      DATAPATH_IxALUOUT_Data1_14_port, DATAPATH_IxALUOUT_Data1_15_port, 
      DATAPATH_IxALUOUT_Data1_16_port, DATAPATH_IxALUOUT_Data1_17_port, 
      DATAPATH_IxALUOUT_Data1_18_port, DATAPATH_IxALUOUT_Data1_19_port, 
      DATAPATH_IxALUOUT_Data1_20_port, DATAPATH_IxALUOUT_Data1_21_port, 
      DATAPATH_IxALUOUT_Data1_22_port, DATAPATH_IxALUOUT_Data1_23_port, 
      DATAPATH_IxALUOUT_Data1_24_port, DATAPATH_IxALUOUT_Data1_25_port, 
      DATAPATH_IxALUOUT_Data1_26_port, DATAPATH_IxALUOUT_Data1_27_port, 
      DATAPATH_IxALUOUT_Data1_28_port, DATAPATH_IxALUOUT_Data1_29_port, 
      DATAPATH_IxALUOUT_Data1_30_port, DATAPATH_IxALUOUT_Data1_31_port, 
      DATAPATH_IxLMD_DATA_0_port, DATAPATH_IxLMD_DATA_1_port, 
      DATAPATH_IxLMD_DATA_2_port, DATAPATH_IxLMD_DATA_3_port, 
      DATAPATH_IxLMD_DATA_4_port, DATAPATH_IxLMD_DATA_5_port, 
      DATAPATH_IxLMD_DATA_6_port, DATAPATH_IxLMD_DATA_7_port, 
      DATAPATH_IxLMD_DATA_8_port, DATAPATH_IxLMD_DATA_9_port, 
      DATAPATH_IxLMD_DATA_10_port, DATAPATH_IxLMD_DATA_11_port, 
      DATAPATH_IxLMD_DATA_12_port, DATAPATH_IxLMD_DATA_13_port, 
      DATAPATH_IxLMD_DATA_14_port, DATAPATH_IxLMD_DATA_15_port, 
      DATAPATH_IxLMD_DATA_16_port, DATAPATH_IxLMD_DATA_17_port, 
      DATAPATH_IxLMD_DATA_18_port, DATAPATH_IxLMD_DATA_19_port, 
      DATAPATH_IxLMD_DATA_20_port, DATAPATH_IxLMD_DATA_21_port, 
      DATAPATH_IxLMD_DATA_22_port, DATAPATH_IxLMD_DATA_23_port, 
      DATAPATH_IxLMD_DATA_24_port, DATAPATH_IxLMD_DATA_25_port, 
      DATAPATH_IxLMD_DATA_26_port, DATAPATH_IxLMD_DATA_27_port, 
      DATAPATH_IxLMD_DATA_28_port, DATAPATH_IxLMD_DATA_29_port, 
      DATAPATH_IxLMD_DATA_30_port, DATAPATH_IxLMD_DATA_31_port, 
      DATAPATH_IxWR_ADD_MEM_fu_0_port, DATAPATH_IxWR_ADD_MEM_fu_1_port, 
      DATAPATH_IxWR_ADD_MEM_fu_2_port, DATAPATH_IxWR_ADD_MEM_fu_3_port, 
      DATAPATH_IxWR_ADD_MEM_fu_4_port, DATAPATH_IxPC4_0_port, 
      DATAPATH_IxPC4_1_port, DATAPATH_IxINSTR_7_port, DATAPATH_IxINSTR_8_port, 
      DATAPATH_IxINSTR_9_port, DATAPATH_IxINSTR_10_port, 
      DATAPATH_IxINSTR_11_port, DATAPATH_IxSecond_stxWRADD_d1_0_port, 
      DATAPATH_IxSecond_stxWRADD_d1_1_port, 
      DATAPATH_IxSecond_stxWRADD_d1_2_port, 
      DATAPATH_IxSecond_stxWRADD_d1_3_port, 
      DATAPATH_IxSecond_stxWRADD_d1_4_port, 
      DATAPATH_IxSecond_stximm_extended_0_port, 
      DATAPATH_IxSecond_stximm_extended_1_port, 
      DATAPATH_IxSecond_stximm_extended_2_port, 
      DATAPATH_IxSecond_stximm_extended_3_port, 
      DATAPATH_IxSecond_stximm_extended_4_port, 
      DATAPATH_IxSecond_stximm_extended_12_port, 
      DATAPATH_IxSecond_stximm_extended_13_port, 
      DATAPATH_IxSecond_stximm_extended_14_port, 
      DATAPATH_IxSecond_stximm_extended_15_port, 
      DATAPATH_IxSecond_stximm_extended_16_port, 
      DATAPATH_IxSecond_stximm_extended_17_port, 
      DATAPATH_IxSecond_stximm_extended_18_port, 
      DATAPATH_IxSecond_stximm_extended_19_port, 
      DATAPATH_IxSecond_stximm_extended_20_port, 
      DATAPATH_IxSecond_stximm_extended_21_port, 
      DATAPATH_IxSecond_stximm_extended_22_port, 
      DATAPATH_IxSecond_stximm_extended_23_port, 
      DATAPATH_IxSecond_stximm_extended_24_port, 
      DATAPATH_IxSecond_stximm_extended_25_port, 
      DATAPATH_IxSecond_stximm_extended_26_port, 
      DATAPATH_IxSecond_stximm_extended_27_port, 
      DATAPATH_IxSecond_stximm_extended_28_port, 
      DATAPATH_IxSecond_stximm_extended_29_port, 
      DATAPATH_IxSecond_stximm_extended_30_port, 
      DATAPATH_IxSecond_stximm_extended_31_port, 
      DATAPATH_IxSecond_stxBR_target_2_port, 
      DATAPATH_IxSecond_stxBR_target_6_port, 
      DATAPATH_IxSecond_stxBR_target_8_port, 
      DATAPATH_IxSecond_stxBR_target_10_port, 
      DATAPATH_IxSecond_stxBR_target_12_port, 
      DATAPATH_IxSecond_stxBR_target_14_port, 
      DATAPATH_IxSecond_stxBR_target_18_port, 
      DATAPATH_IxSecond_stxjump_target_0_port, 
      DATAPATH_IxSecond_stxjump_target_3_port, 
      DATAPATH_IxSecond_stxjump_target_5_port, 
      DATAPATH_IxSecond_stxjump_target_6_port, 
      DATAPATH_IxSecond_stxjump_target_7_port, 
      DATAPATH_IxSecond_stxjump_target_10_port, 
      DATAPATH_IxSecond_stxjump_target_11_port, 
      DATAPATH_IxSecond_stxjump_target_12_port, 
      DATAPATH_IxSecond_stxjump_target_14_port, 
      DATAPATH_IxSecond_stxjump_target_16_port, 
      DATAPATH_IxSecond_stxjump_target_17_port, 
      DATAPATH_IxSecond_stxjump_target_18_port, 
      DATAPATH_IxSecond_stxjump_target_21_port, 
      DATAPATH_IxSecond_stxjump_target_22_port, 
      DATAPATH_IxSecond_stxjump_target_23_port, 
      DATAPATH_IxSecond_stxjump_target_25_port, 
      DATAPATH_IxSecond_stxjump_target_26_port, 
      DATAPATH_IxSecond_stxjump_target_27_port, 
      DATAPATH_IxSecond_stxjump_target_30_port, 
      DATAPATH_IxSecond_stxjump_target_31_port, 
      DATAPATH_IxThird_stxALU_out_i_0_port, 
      DATAPATH_IxThird_stxALU_out_i_1_port, 
      DATAPATH_IxThird_stxALU_out_i_2_port, 
      DATAPATH_IxThird_stxALU_out_i_3_port, 
      DATAPATH_IxThird_stxALU_out_i_4_port, 
      DATAPATH_IxThird_stxALU_out_i_5_port, 
      DATAPATH_IxThird_stxALU_out_i_6_port, 
      DATAPATH_IxThird_stxALU_out_i_7_port, 
      DATAPATH_IxThird_stxALU_out_i_8_port, 
      DATAPATH_IxThird_stxALU_out_i_9_port, 
      DATAPATH_IxThird_stxALU_out_i_10_port, 
      DATAPATH_IxThird_stxALU_out_i_11_port, 
      DATAPATH_IxThird_stxALU_out_i_12_port, 
      DATAPATH_IxThird_stxALU_out_i_13_port, 
      DATAPATH_IxThird_stxALU_out_i_14_port, 
      DATAPATH_IxThird_stxALU_out_i_15_port, 
      DATAPATH_IxThird_stxALU_out_i_16_port, 
      DATAPATH_IxThird_stxALU_out_i_17_port, 
      DATAPATH_IxThird_stxALU_out_i_18_port, 
      DATAPATH_IxThird_stxALU_out_i_19_port, 
      DATAPATH_IxThird_stxALU_out_i_20_port, 
      DATAPATH_IxThird_stxALU_out_i_21_port, 
      DATAPATH_IxThird_stxALU_out_i_22_port, 
      DATAPATH_IxThird_stxALU_out_i_23_port, 
      DATAPATH_IxThird_stxALU_out_i_24_port, 
      DATAPATH_IxThird_stxALU_out_i_25_port, 
      DATAPATH_IxThird_stxALU_out_i_26_port, 
      DATAPATH_IxThird_stxALU_out_i_27_port, 
      DATAPATH_IxThird_stxALU_out_i_28_port, 
      DATAPATH_IxThird_stxALU_out_i_29_port, 
      DATAPATH_IxThird_stxALU_out_i_30_port, 
      DATAPATH_IxThird_stxALU_out_i_31_port, DATAPATH_IxThird_stxALU_IN2_0_port
      , DATAPATH_IxThird_stxALU_IN2_1_port, DATAPATH_IxThird_stxALU_IN2_2_port,
      DATAPATH_IxThird_stxALU_IN2_3_port, DATAPATH_IxThird_stxALU_IN2_4_port, 
      DATAPATH_IxThird_stxALU_IN2_5_port, DATAPATH_IxThird_stxALU_IN1_0_port, 
      DATAPATH_IxThird_stxALU_IN1_1_port, DATAPATH_IxThird_stxALU_IN1_2_port, 
      DATAPATH_IxThird_stxALU_IN1_3_port, DATAPATH_IxThird_stxALU_IN1_4_port, 
      DATAPATH_IxThird_stxALU_IN1_5_port, DATAPATH_IxThird_stxALU_IN1_6_port, 
      DATAPATH_IxThird_stxALU_IN1_7_port, DATAPATH_IxThird_stxALU_IN1_8_port, 
      DATAPATH_IxThird_stxALU_IN1_9_port, DATAPATH_IxThird_stxALU_IN1_10_port, 
      DATAPATH_IxThird_stxALU_IN1_11_port, DATAPATH_IxThird_stxALU_IN1_12_port,
      DATAPATH_IxThird_stxALU_IN1_13_port, DATAPATH_IxThird_stxALU_IN1_14_port,
      DATAPATH_IxThird_stxALU_IN1_15_port, DATAPATH_IxThird_stxALU_IN1_16_port,
      DATAPATH_IxThird_stxALU_IN1_17_port, DATAPATH_IxThird_stxALU_IN1_18_port,
      DATAPATH_IxThird_stxALU_IN1_19_port, DATAPATH_IxThird_stxALU_IN1_20_port,
      DATAPATH_IxThird_stxALU_IN1_21_port, DATAPATH_IxThird_stxALU_IN1_22_port,
      DATAPATH_IxThird_stxALU_IN1_23_port, DATAPATH_IxThird_stxALU_IN1_24_port,
      DATAPATH_IxThird_stxALU_IN1_25_port, DATAPATH_IxThird_stxALU_IN1_26_port,
      DATAPATH_IxThird_stxALU_IN1_27_port, DATAPATH_IxThird_stxALU_IN1_28_port,
      DATAPATH_IxThird_stxALU_IN1_29_port, DATAPATH_IxThird_stxALU_IN1_30_port,
      DATAPATH_IxThird_stxALU1xN222, DATAPATH_IxThird_stxALU1xN221, 
      DATAPATH_IxThird_stxALU1xN220, DATAPATH_IxThird_stxALU1xN219, 
      DATAPATH_IxThird_stxALU1xN218, DATAPATH_IxThird_stxALU1xN217, 
      DATAPATH_IxThird_stxALU1xN216, DATAPATH_IxThird_stxALU1xN215, 
      DATAPATH_IxThird_stxALU1xN214, DATAPATH_IxThird_stxALU1xN213, 
      DATAPATH_IxThird_stxALU1xN212, DATAPATH_IxThird_stxALU1xN211, 
      DATAPATH_IxThird_stxALU1xN210, DATAPATH_IxThird_stxALU1xN209, 
      DATAPATH_IxThird_stxALU1xN208, DATAPATH_IxThird_stxALU1xN207, 
      DATAPATH_IxThird_stxALU1xN206, DATAPATH_IxThird_stxALU1xN205, 
      DATAPATH_IxThird_stxALU1xN204, DATAPATH_IxThird_stxALU1xN203, 
      DATAPATH_IxThird_stxALU1xN202, DATAPATH_IxThird_stxALU1xN201, 
      DATAPATH_IxThird_stxALU1xN200, DATAPATH_IxThird_stxALU1xN199, 
      DATAPATH_IxThird_stxALU1xN198, DATAPATH_IxThird_stxALU1xN197, 
      DATAPATH_IxThird_stxALU1xN196, DATAPATH_IxThird_stxALU1xN195, 
      DATAPATH_IxThird_stxALU1xN194, DATAPATH_IxThird_stxALU1xN193, 
      DATAPATH_IxThird_stxALU1xN192, DATAPATH_IxThird_stxALU1xN191, n22, n23, 
      n25, n26, n27, n28, n29, n32, n33, n35, n36, n37, n38, n43, n46, n47, n48
      , n49, n54, n91, n92, n96, n97, n99, n101, n103, n105, n106, n108, n109, 
      n110, n111, n112, n113, n115, n118, n119, n120, n122, n124, n126, n129, 
      n130, n132, n134, n135, n137, n139, n141, n143, n144, n145, n146, n148, 
      n150, n152, n154, n156, n158, n159, n160, n161, n162, n164, n165, n167, 
      n168, n169, n171, n172, n174, n175, n177, n179, n180, n181, n182, n183, 
      n185, n187, n188, n189, n190, n191, n192, n194, n196, n197, n198, n200, 
      n201, n203, n205, n206, n207, n209, n211, n212, n213, n214, n216, n217, 
      n218, n219, n221, n222, n223, n224, n226, n228, n229, n231, n232, n233, 
      n234, n236, n237, n238, n239, n241, n242, n243, n244, n246, n248, n250, 
      n251, n253, n254, n255, n256, n258, n260, n261, n262, n265, n266, n267, 
      n268, n269, n270, n271, n273, n275, n278, n279, n280, n282, n283, n284, 
      n285, n286, n289, n291, n292, n294, n296, n298, n299, n326, n328, n330, 
      n331, n333, n334, n335, n336, n337, n338, n340, n344, n345, n346, n347, 
      n348, n349, n351, n352, n353, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n367, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n382, n383, n384, n385, n386, n387, n388, 
      n390, n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n411, n412, n413, n416, n418, n419, n420, 
      n421, n422, n423, n425, n426, n427, n428, n429, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n446, n447, 
      n449, n450, n451, n452, n453, n454, n455, n457, n459, n460, n461, n463, 
      n464, n465, n467, n468, n469, n470, n471, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n483, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n495, n496, n497, n498, n500, n501, n502, n503, n504, n505, 
      n507, n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520, 
      n522, n523, n524, n525, n526, n527, n528, n529, n530, n532, n534, n535, 
      n536, n537, n538, n539, n540, n541, n543, n544, n545, n546, n548, n549, 
      n550, n551, n552, n553, n555, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n567, n568, n569, n570, n571, n572, n574, n575, n576, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n590, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n605, n607, 
      n608, n609, n610, n611, n613, n615, n616, n617, n618, n619, n620, n622, 
      n623, n624, n625, n626, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n638, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n652, n653, n654, n655, n656, n657, n658, n660, n661, n662, n663, 
      n664, n665, n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n682, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n695, n696, n698, n699, n700, n702, n703, n705, n706, n707, 
      n708, n709, n710, n712, n713, n715, n716, n717, n718, n719, n722, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n737, n738, 
      n739, n740, n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, 
      n753, n754, n755, n757, n758, n759, n760, n762, n763, n765, n766, n767, 
      n768, n769, n770, n771, n773, n774, n775, n776, n778, n779, n780, n781, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n794, n795, 
      n797, n798, n799, n800, n801, n803, n804, n805, n806, n807, n808, n809, 
      n811, n812, n813, n814, n815, n817, n818, n819, n820, n821, n822, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n843, n844, n845, n846, n847, n848, n849, 
      n850, n851, n852, n853, n854, n855, n857, n858, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n876, 
      n877, n878, n879, n882, n884, n885, n886, n887, n889, n890, n894, n896, 
      n897, n898, n899, n900, n901, n903, n904, n905, n906, n907, n909, n910, 
      n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, 
      n924, n925, n927, n929, n930, n931, n932, n933, n934, n936, n938, n939, 
      n940, n941, n942, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n956, n958, n959, n961, n962, n963, n965, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n976, n977, n979, n980, n981, n982, 
      n983, n985, n986, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088, 
      n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1111, 
      n1113, n1114, n1115, n1116, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1137, n1138, n1139, n1140, n1141, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
      n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
      n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1241, n1244, 
      n1248, n1257, n1274, n1275, n1276, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1291, n1292, n1296, n1298, n1299, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, RF_WR_DATAx0x, RF_WR_DATAx1x, RF_WR_DATAx2x, RF_WR_DATAx3x,
      RF_WR_DATAx4x, RF_WR_DATAx5x, RF_WR_DATAx6x, RF_WR_DATAx7x, RF_WR_DATAx8x
      , RF_WR_DATAx9x, RF_WR_DATAx10x, RF_WR_DATAx11x, RF_WR_DATAx12x, 
      RF_WR_DATAx13x, RF_WR_DATAx14x, RF_WR_DATAx15x, RF_WR_DATAx16x, 
      RF_WR_DATAx17x, RF_WR_DATAx18x, RF_WR_DATAx19x, RF_WR_DATAx20x, 
      RF_WR_DATAx21x, RF_WR_DATAx22x, RF_WR_DATAx23x, RF_WR_DATAx24x, 
      RF_WR_DATAx25x, RF_WR_DATAx26x, RF_WR_DATAx27x, RF_WR_DATAx28x, 
      RF_WR_DATAx29x, RF_WR_DATAx30x, RF_WR_DATAx31x, n1961, n1962, n1963, 
      n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, 
      n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, 
      n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
      n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, 
      n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
      n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
      n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, 
      n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
      n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, 
      n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, 
      n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
      n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263 : std_logic;

begin
   IRAM_ADD <= ( IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, DATAPATH_IxPC4_1_port,
      DATAPATH_IxPC4_0_port );
   RF_RD1_ADD <= ( RF_RD1_ADD_4_port, RF_RD1_ADD_3_port, RF_RD1_ADD_2_port, 
      RF_RD1_ADD_1_port, RF_RD1_ADD_0_port );
   RF_RD2_ADD <= ( RF_RD2_ADD_4_port, RF_RD2_ADD_3_port, RF_RD2_ADD_2_port, 
      RF_RD2_ADD_1_port, RF_RD2_ADD_0_port );
   RF_WR_DATA <= ( RF_WR_DATAx31x, RF_WR_DATAx30x, RF_WR_DATAx29x, 
      RF_WR_DATAx28x, RF_WR_DATAx27x, RF_WR_DATAx26x, RF_WR_DATAx25x, 
      RF_WR_DATAx24x, RF_WR_DATAx23x, RF_WR_DATAx22x, RF_WR_DATAx21x, 
      RF_WR_DATAx20x, RF_WR_DATAx19x, RF_WR_DATAx18x, RF_WR_DATAx17x, 
      RF_WR_DATAx16x, RF_WR_DATAx15x, RF_WR_DATAx14x, RF_WR_DATAx13x, 
      RF_WR_DATAx12x, RF_WR_DATAx11x, RF_WR_DATAx10x, RF_WR_DATAx9x, 
      RF_WR_DATAx8x, RF_WR_DATAx7x, RF_WR_DATAx6x, RF_WR_DATAx5x, RF_WR_DATAx4x
      , RF_WR_DATAx3x, RF_WR_DATAx2x, RF_WR_DATAx1x, RF_WR_DATAx0x );
   DRAM_ADD <= ( DRAM_ADD_31_port, DRAM_ADD_30_port, DRAM_ADD_29_port, 
      DRAM_ADD_28_port, DRAM_ADD_27_port, DRAM_ADD_26_port, DRAM_ADD_25_port, 
      DRAM_ADD_24_port, DRAM_ADD_23_port, DRAM_ADD_22_port, DRAM_ADD_21_port, 
      DRAM_ADD_20_port, DRAM_ADD_19_port, DRAM_ADD_18_port, DRAM_ADD_17_port, 
      DRAM_ADD_16_port, DRAM_ADD_15_port, DRAM_ADD_14_port, DRAM_ADD_13_port, 
      DRAM_ADD_12_port, DRAM_ADD_11_port, DRAM_ADD_10_port, DRAM_ADD_9_port, 
      DRAM_ADD_8_port, DRAM_ADD_7_port, DRAM_ADD_6_port, DRAM_ADD_5_port, 
      DRAM_ADD_4_port, DRAM_ADD_3_port, DRAM_ADD_2_port, DRAM_ADD_1_port, 
      DRAM_ADD_0_port );
   
   CU_IxaluOpcode2_regx0x : DFF_X1 port map( D => n1289, CK => Clk, Q => n1623,
                           QN => n1276);
   CU_IxaluOpcode2_regx1x : DFF_X1 port map( D => n1288, CK => Clk, Q => n_1000
                           , QN => n1275);
   CU_IxaluOpcode2_regx2x : DFF_X1 port map( D => n1287, CK => Clk, Q => n_1001
                           , QN => n1274);
   CU_IxaluOpcode3_regx0x : DFF_X1 port map( D => n1286, CK => Clk, Q => n_1002
                           , QN => n1335);
   CU_IxaluOpcode3_regx1x : DFF_X1 port map( D => n1285, CK => Clk, Q => n1591,
                           QN => n1336);
   CU_IxaluOpcode3_regx2x : DFF_X1 port map( D => n1284, CK => Clk, Q => n1613,
                           QN => n1337);
   DATAPATH_IxThird_stxB_FORWARD_out_regx0x : DFF_X1 port map( D => 
                           RF_RD2_DATA(0), CK => Clk, Q => DRAM_DIN(0), QN => 
                           n_1003);
   DATAPATH_IxThird_stxB_FORWARD_out_regx1x : DFF_X1 port map( D => 
                           RF_RD2_DATA(1), CK => Clk, Q => DRAM_DIN(1), QN => 
                           n_1004);
   DATAPATH_IxThird_stxB_FORWARD_out_regx2x : DFF_X1 port map( D => 
                           RF_RD2_DATA(2), CK => Clk, Q => DRAM_DIN(2), QN => 
                           n_1005);
   DATAPATH_IxThird_stxB_FORWARD_out_regx3x : DFF_X1 port map( D => 
                           RF_RD2_DATA(3), CK => Clk, Q => DRAM_DIN(3), QN => 
                           n_1006);
   DATAPATH_IxThird_stxB_FORWARD_out_regx4x : DFF_X1 port map( D => 
                           RF_RD2_DATA(4), CK => Clk, Q => DRAM_DIN(4), QN => 
                           n_1007);
   DATAPATH_IxThird_stxB_FORWARD_out_regx5x : DFF_X1 port map( D => 
                           RF_RD2_DATA(5), CK => Clk, Q => DRAM_DIN(5), QN => 
                           n_1008);
   DATAPATH_IxThird_stxB_FORWARD_out_regx6x : DFF_X1 port map( D => 
                           RF_RD2_DATA(6), CK => Clk, Q => DRAM_DIN(6), QN => 
                           n_1009);
   DATAPATH_IxThird_stxB_FORWARD_out_regx7x : DFF_X1 port map( D => 
                           RF_RD2_DATA(7), CK => Clk, Q => DRAM_DIN(7), QN => 
                           n_1010);
   DATAPATH_IxThird_stxB_FORWARD_out_regx8x : DFF_X1 port map( D => 
                           RF_RD2_DATA(8), CK => Clk, Q => DRAM_DIN(8), QN => 
                           n_1011);
   DATAPATH_IxThird_stxB_FORWARD_out_regx9x : DFF_X1 port map( D => 
                           RF_RD2_DATA(9), CK => Clk, Q => DRAM_DIN(9), QN => 
                           n_1012);
   DATAPATH_IxThird_stxB_FORWARD_out_regx10x : DFF_X1 port map( D => 
                           RF_RD2_DATA(10), CK => Clk, Q => DRAM_DIN(10), QN =>
                           n_1013);
   DATAPATH_IxThird_stxB_FORWARD_out_regx11x : DFF_X1 port map( D => 
                           RF_RD2_DATA(11), CK => Clk, Q => DRAM_DIN(11), QN =>
                           n_1014);
   DATAPATH_IxThird_stxB_FORWARD_out_regx12x : DFF_X1 port map( D => 
                           RF_RD2_DATA(12), CK => Clk, Q => DRAM_DIN(12), QN =>
                           n_1015);
   DATAPATH_IxThird_stxB_FORWARD_out_regx13x : DFF_X1 port map( D => 
                           RF_RD2_DATA(13), CK => Clk, Q => DRAM_DIN(13), QN =>
                           n_1016);
   DATAPATH_IxThird_stxB_FORWARD_out_regx14x : DFF_X1 port map( D => 
                           RF_RD2_DATA(14), CK => Clk, Q => DRAM_DIN(14), QN =>
                           n_1017);
   DATAPATH_IxThird_stxB_FORWARD_out_regx15x : DFF_X1 port map( D => 
                           RF_RD2_DATA(15), CK => Clk, Q => DRAM_DIN(15), QN =>
                           n_1018);
   DATAPATH_IxThird_stxB_FORWARD_out_regx16x : DFF_X1 port map( D => 
                           RF_RD2_DATA(16), CK => Clk, Q => DRAM_DIN(16), QN =>
                           n_1019);
   DATAPATH_IxThird_stxB_FORWARD_out_regx17x : DFF_X1 port map( D => 
                           RF_RD2_DATA(17), CK => Clk, Q => DRAM_DIN(17), QN =>
                           n_1020);
   DATAPATH_IxThird_stxB_FORWARD_out_regx18x : DFF_X1 port map( D => 
                           RF_RD2_DATA(18), CK => Clk, Q => DRAM_DIN(18), QN =>
                           n_1021);
   DATAPATH_IxThird_stxB_FORWARD_out_regx19x : DFF_X1 port map( D => 
                           RF_RD2_DATA(19), CK => Clk, Q => DRAM_DIN(19), QN =>
                           n_1022);
   DATAPATH_IxThird_stxB_FORWARD_out_regx20x : DFF_X1 port map( D => 
                           RF_RD2_DATA(20), CK => Clk, Q => DRAM_DIN(20), QN =>
                           n_1023);
   DATAPATH_IxThird_stxB_FORWARD_out_regx21x : DFF_X1 port map( D => 
                           RF_RD2_DATA(21), CK => Clk, Q => DRAM_DIN(21), QN =>
                           n_1024);
   DATAPATH_IxThird_stxB_FORWARD_out_regx22x : DFF_X1 port map( D => 
                           RF_RD2_DATA(22), CK => Clk, Q => DRAM_DIN(22), QN =>
                           n_1025);
   DATAPATH_IxThird_stxB_FORWARD_out_regx23x : DFF_X1 port map( D => 
                           RF_RD2_DATA(23), CK => Clk, Q => DRAM_DIN(23), QN =>
                           n_1026);
   DATAPATH_IxThird_stxB_FORWARD_out_regx24x : DFF_X1 port map( D => 
                           RF_RD2_DATA(24), CK => Clk, Q => DRAM_DIN(24), QN =>
                           n_1027);
   DATAPATH_IxThird_stxB_FORWARD_out_regx25x : DFF_X1 port map( D => 
                           RF_RD2_DATA(25), CK => Clk, Q => DRAM_DIN(25), QN =>
                           n_1028);
   DATAPATH_IxThird_stxB_FORWARD_out_regx26x : DFF_X1 port map( D => 
                           RF_RD2_DATA(26), CK => Clk, Q => DRAM_DIN(26), QN =>
                           n_1029);
   DATAPATH_IxThird_stxB_FORWARD_out_regx27x : DFF_X1 port map( D => 
                           RF_RD2_DATA(27), CK => Clk, Q => DRAM_DIN(27), QN =>
                           n_1030);
   DATAPATH_IxThird_stxB_FORWARD_out_regx28x : DFF_X1 port map( D => 
                           RF_RD2_DATA(28), CK => Clk, Q => DRAM_DIN(28), QN =>
                           n_1031);
   DATAPATH_IxThird_stxB_FORWARD_out_regx29x : DFF_X1 port map( D => 
                           RF_RD2_DATA(29), CK => Clk, Q => DRAM_DIN(29), QN =>
                           n_1032);
   DATAPATH_IxThird_stxB_FORWARD_out_regx30x : DFF_X1 port map( D => 
                           RF_RD2_DATA(30), CK => Clk, Q => DRAM_DIN(30), QN =>
                           n_1033);
   DATAPATH_IxThird_stxB_FORWARD_out_regx31x : DFF_X1 port map( D => 
                           RF_RD2_DATA(31), CK => Clk, Q => DRAM_DIN(31), QN =>
                           n_1034);
   DATAPATH_IxFourth_stxLMD_out_regx0x : DFF_X1 port map( D => DRAM_DOUT(0), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_0_port, QN => 
                           n_1035);
   DATAPATH_IxFourth_stxLMD_out_regx1x : DFF_X1 port map( D => DRAM_DOUT(1), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_1_port, QN => 
                           n_1036);
   DATAPATH_IxFourth_stxLMD_out_regx2x : DFF_X1 port map( D => DRAM_DOUT(2), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_2_port, QN => 
                           n_1037);
   DATAPATH_IxFourth_stxLMD_out_regx3x : DFF_X1 port map( D => DRAM_DOUT(3), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_3_port, QN => 
                           n_1038);
   DATAPATH_IxFourth_stxLMD_out_regx4x : DFF_X1 port map( D => DRAM_DOUT(4), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_4_port, QN => 
                           n_1039);
   DATAPATH_IxFourth_stxLMD_out_regx5x : DFF_X1 port map( D => DRAM_DOUT(5), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_5_port, QN => 
                           n_1040);
   DATAPATH_IxFourth_stxLMD_out_regx6x : DFF_X1 port map( D => DRAM_DOUT(6), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_6_port, QN => 
                           n_1041);
   DATAPATH_IxFourth_stxLMD_out_regx7x : DFF_X1 port map( D => DRAM_DOUT(7), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_7_port, QN => 
                           n_1042);
   DATAPATH_IxFourth_stxLMD_out_regx8x : DFF_X1 port map( D => DRAM_DOUT(8), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_8_port, QN => 
                           n_1043);
   DATAPATH_IxFourth_stxLMD_out_regx9x : DFF_X1 port map( D => DRAM_DOUT(9), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_9_port, QN => 
                           n_1044);
   DATAPATH_IxFourth_stxLMD_out_regx10x : DFF_X1 port map( D => DRAM_DOUT(10), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_10_port, QN => 
                           n_1045);
   DATAPATH_IxFourth_stxLMD_out_regx11x : DFF_X1 port map( D => DRAM_DOUT(11), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_11_port, QN => 
                           n_1046);
   DATAPATH_IxFourth_stxLMD_out_regx12x : DFF_X1 port map( D => DRAM_DOUT(12), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_12_port, QN => 
                           n_1047);
   DATAPATH_IxFourth_stxLMD_out_regx13x : DFF_X1 port map( D => DRAM_DOUT(13), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_13_port, QN => 
                           n_1048);
   DATAPATH_IxFourth_stxLMD_out_regx14x : DFF_X1 port map( D => DRAM_DOUT(14), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_14_port, QN => 
                           n_1049);
   DATAPATH_IxFourth_stxLMD_out_regx15x : DFF_X1 port map( D => DRAM_DOUT(15), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_15_port, QN => 
                           n_1050);
   DATAPATH_IxFourth_stxLMD_out_regx16x : DFF_X1 port map( D => DRAM_DOUT(16), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_16_port, QN => 
                           n_1051);
   DATAPATH_IxFourth_stxLMD_out_regx17x : DFF_X1 port map( D => DRAM_DOUT(17), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_17_port, QN => 
                           n_1052);
   DATAPATH_IxFourth_stxLMD_out_regx18x : DFF_X1 port map( D => DRAM_DOUT(18), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_18_port, QN => 
                           n_1053);
   DATAPATH_IxFourth_stxLMD_out_regx19x : DFF_X1 port map( D => DRAM_DOUT(19), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_19_port, QN => 
                           n_1054);
   DATAPATH_IxFourth_stxLMD_out_regx20x : DFF_X1 port map( D => DRAM_DOUT(20), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_20_port, QN => 
                           n_1055);
   DATAPATH_IxFourth_stxLMD_out_regx21x : DFF_X1 port map( D => DRAM_DOUT(21), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_21_port, QN => 
                           n_1056);
   DATAPATH_IxFourth_stxLMD_out_regx22x : DFF_X1 port map( D => DRAM_DOUT(22), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_22_port, QN => 
                           n_1057);
   DATAPATH_IxFourth_stxLMD_out_regx23x : DFF_X1 port map( D => DRAM_DOUT(23), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_23_port, QN => 
                           n_1058);
   DATAPATH_IxFourth_stxLMD_out_regx24x : DFF_X1 port map( D => DRAM_DOUT(24), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_24_port, QN => 
                           n_1059);
   DATAPATH_IxFourth_stxLMD_out_regx25x : DFF_X1 port map( D => DRAM_DOUT(25), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_25_port, QN => 
                           n_1060);
   DATAPATH_IxFourth_stxLMD_out_regx26x : DFF_X1 port map( D => DRAM_DOUT(26), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_26_port, QN => 
                           n_1061);
   DATAPATH_IxFourth_stxLMD_out_regx27x : DFF_X1 port map( D => DRAM_DOUT(27), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_27_port, QN => 
                           n_1062);
   DATAPATH_IxFourth_stxLMD_out_regx28x : DFF_X1 port map( D => DRAM_DOUT(28), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_28_port, QN => 
                           n_1063);
   DATAPATH_IxFourth_stxLMD_out_regx29x : DFF_X1 port map( D => DRAM_DOUT(29), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_29_port, QN => 
                           n_1064);
   DATAPATH_IxFourth_stxLMD_out_regx30x : DFF_X1 port map( D => DRAM_DOUT(30), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_30_port, QN => 
                           n_1065);
   DATAPATH_IxFourth_stxLMD_out_regx31x : DFF_X1 port map( D => DRAM_DOUT(31), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_31_port, QN => 
                           n_1066);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_0_port, CK => Clk, Q 
                           => DRAM_ADD_0_port, QN => n1419);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx0x : DFF_X1 port map( D => 
                           DRAM_ADD_0_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_0_port, QN => n_1067);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx10x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_10_port, CK => Clk, Q 
                           => DRAM_ADD_10_port, QN => n1429);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx10x : DFF_X1 port map( D => 
                           DRAM_ADD_10_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_10_port, QN => n_1068);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_16_port, CK => Clk, Q 
                           => DRAM_ADD_16_port, QN => n1435);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx16x : DFF_X1 port map( D => 
                           DRAM_ADD_16_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_16_port, QN => n_1069);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_17_port, CK => Clk, Q 
                           => DRAM_ADD_17_port, QN => n1436);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx17x : DFF_X1 port map( D => 
                           DRAM_ADD_17_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_17_port, QN => n_1070);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_18_port, CK => Clk, Q 
                           => DRAM_ADD_18_port, QN => n1437);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx18x : DFF_X1 port map( D => 
                           DRAM_ADD_18_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_18_port, QN => n_1071);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_25_port, CK => Clk, Q 
                           => DRAM_ADD_25_port, QN => n1444);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx25x : DFF_X1 port map( D => 
                           DRAM_ADD_25_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_25_port, QN => n_1072);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_26_port, CK => Clk, Q 
                           => DRAM_ADD_26_port, QN => n1445);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx26x : DFF_X1 port map( D => 
                           DRAM_ADD_26_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_26_port, QN => n_1073);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_31_port, CK => Clk, Q 
                           => DRAM_ADD_31_port, QN => n1450);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx31x : DFF_X1 port map( D => 
                           DRAM_ADD_31_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_31_port, QN => n_1074);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx31x : DFF_X1 port map( D => n1548, CK 
                           => Clk, Q => n1621, QN => n1386);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx30x : DFF_X1 port map( D => n1549, CK 
                           => Clk, Q => n_1075, QN => n1385);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx29x : DFF_X1 port map( D => n1550, CK 
                           => Clk, Q => n_1076, QN => n1624);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx28x : DFF_X1 port map( D => n1551, CK 
                           => Clk, Q => n_1077, QN => n1384);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx27x : DFF_X1 port map( D => n1552, CK 
                           => Clk, Q => n_1078, QN => n1383);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx26x : DFF_X1 port map( D => n1553, CK 
                           => Clk, Q => n_1079, QN => n1382);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx25x : DFF_X1 port map( D => n1554, CK 
                           => Clk, Q => n_1080, QN => n1381);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx24x : DFF_X1 port map( D => n1555, CK 
                           => Clk, Q => RF_RD2_ADD_4_port, QN => n1380);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx4x : DFF_X1 port map( D => 
                           RF_RD2_ADD_4_port, CK => Clk, Q => n_1081, QN => 
                           n1154);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx23x : DFF_X1 port map( D => n1556, CK 
                           => Clk, Q => RF_RD2_ADD_3_port, QN => n1379);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx3x : DFF_X1 port map( D => 
                           RF_RD2_ADD_3_port, CK => Clk, Q => n_1082, QN => 
                           n1156);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx22x : DFF_X1 port map( D => n1557, CK 
                           => Clk, Q => RF_RD2_ADD_2_port, QN => n1378);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx2x : DFF_X1 port map( D => 
                           RF_RD2_ADD_2_port, CK => Clk, Q => n_1083, QN => 
                           n1153);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx21x : DFF_X1 port map( D => n1558, CK 
                           => Clk, Q => RF_RD2_ADD_1_port, QN => n1377);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx1x : DFF_X1 port map( D => 
                           RF_RD2_ADD_1_port, CK => Clk, Q => n_1084, QN => 
                           n1155);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx20x : DFF_X1 port map( D => n1559, CK 
                           => Clk, Q => RF_RD2_ADD_0_port, QN => n1376);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx0x : DFF_X1 port map( D => 
                           RF_RD2_ADD_0_port, CK => Clk, Q => n_1085, QN => 
                           n1152);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx19x : DFF_X1 port map( D => n1560, CK 
                           => Clk, Q => RF_RD1_ADD_4_port, QN => n1375);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx4x : DFF_X1 port map( D => 
                           RF_RD1_ADD_4_port, CK => Clk, Q => n_1086, QN => 
                           n1164);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx18x : DFF_X1 port map( D => n1561, CK 
                           => Clk, Q => RF_RD1_ADD_3_port, QN => n1374);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx3x : DFF_X1 port map( D => 
                           RF_RD1_ADD_3_port, CK => Clk, Q => n_1087, QN => 
                           n1165);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx17x : DFF_X1 port map( D => n1562, CK 
                           => Clk, Q => RF_RD1_ADD_2_port, QN => n1373);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx2x : DFF_X1 port map( D => 
                           RF_RD1_ADD_2_port, CK => Clk, Q => n_1088, QN => 
                           n1163);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx16x : DFF_X1 port map( D => n1563, CK 
                           => Clk, Q => RF_RD1_ADD_1_port, QN => n1372);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx1x : DFF_X1 port map( D => 
                           RF_RD1_ADD_1_port, CK => Clk, Q => n_1089, QN => 
                           n1162);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx15x : DFF_X1 port map( D => n1564, CK 
                           => Clk, Q => RF_RD1_ADD_0_port, QN => n1371);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx0x : DFF_X1 port map( D => 
                           RF_RD1_ADD_0_port, CK => Clk, Q => n_1090, QN => 
                           n1161);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx14x : DFF_X1 port map( D => n1565, CK 
                           => Clk, Q => n1210, QN => n1615);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx13x : DFF_X1 port map( D => n1566, CK 
                           => Clk, Q => n_1091, QN => n1609);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx12x : DFF_X1 port map( D => n1567, CK 
                           => Clk, Q => n_1092, QN => n1608);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx11x : DFF_X1 port map( D => n1568, CK 
                           => Clk, Q => DATAPATH_IxINSTR_11_port, QN => n1370);
   DATAPATH_IxSecond_stxWRADD_d1_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_11_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, QN => n_1093);
   DATAPATH_IxSecond_stxWRADD_d2_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_4_port, QN => n1150);
   DATAPATH_IxSecond_stxWRADD_d3_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_4_port, CK => Clk, Q => 
                           RF_WR_ADD(4), QN => n1158);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx10x : DFF_X1 port map( D => n1569, CK 
                           => Clk, Q => DATAPATH_IxINSTR_10_port, QN => n1369);
   DATAPATH_IxSecond_stxWRADD_d1_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_10_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, QN => n_1094);
   DATAPATH_IxSecond_stxWRADD_d2_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_3_port, QN => n1149);
   DATAPATH_IxSecond_stxWRADD_d3_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_3_port, CK => Clk, Q => 
                           RF_WR_ADD(3), QN => n1160);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx9x : DFF_X1 port map( D => n1570, CK =>
                           Clk, Q => DATAPATH_IxINSTR_9_port, QN => n1368);
   DATAPATH_IxSecond_stxWRADD_d1_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_9_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, QN => n_1095);
   DATAPATH_IxSecond_stxWRADD_d2_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_2_port, QN => n1147);
   DATAPATH_IxSecond_stxWRADD_d3_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_2_port, CK => Clk, Q => 
                           RF_WR_ADD(2), QN => n1146);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx8x : DFF_X1 port map( D => n1571, CK =>
                           Clk, Q => DATAPATH_IxINSTR_8_port, QN => n1367);
   DATAPATH_IxSecond_stxWRADD_d1_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_8_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, QN => n_1096);
   DATAPATH_IxSecond_stxWRADD_d2_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_1_port, QN => n1148);
   DATAPATH_IxSecond_stxWRADD_d3_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_1_port, CK => Clk, Q => 
                           RF_WR_ADD(1), QN => n1159);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx7x : DFF_X1 port map( D => n1572, CK =>
                           Clk, Q => DATAPATH_IxINSTR_7_port, QN => n1366);
   DATAPATH_IxSecond_stxWRADD_d1_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_7_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, QN => n_1097);
   DATAPATH_IxSecond_stxWRADD_d2_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_0_port, QN => n1151);
   DATAPATH_IxSecond_stxWRADD_d3_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_0_port, CK => Clk, Q => 
                           RF_WR_ADD(0), QN => n1145);
   CU_Ixcw2_i_regx12x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1743, Q => CU_Ixcw2_i_12_port, QN => n_1098);
   CU_Ixcw3_regx5x : DFFR_X1 port map( D => CU_Ixcw2_5_port, CK => Clk, RN => 
                           n1744, Q => IMM_SEL_i, QN => n_1099);
   CU_Ixcw3_regx4x : DFFR_X1 port map( D => CU_Ixcw2_4_port, CK => Clk, RN => 
                           n1744, Q => BRANCH_EN_i, QN => n_1100);
   CU_Ixcw3_regx3x : DFFR_X1 port map( D => CU_Ixcw2_3_port, CK => Clk, RN => 
                           n1744, Q => CU_Ixcw3_3_port, QN => n_1101);
   CU_Ixcw4_regx3x : DFFR_X1 port map( D => CU_Ixcw3_3_port, CK => Clk, RN => 
                           n1744, Q => DRAM_WE, QN => n_1102);
   CU_Ixcw3_regx2x : DFFR_X1 port map( D => CU_Ixcw2_2_port, CK => Clk, RN => 
                           n1744, Q => CU_Ixcw3_2_port, QN => n_1103);
   CU_Ixcw4_regx2x : DFFR_X1 port map( D => CU_Ixcw3_2_port, CK => Clk, RN => 
                           n1743, Q => DRAM_RE, QN => n_1104);
   CU_Ixcw3_regx1x : DFFR_X1 port map( D => CU_Ixcw2_1_port, CK => Clk, RN => 
                           n1744, Q => CU_Ixcw3_1_port, QN => n_1105);
   CU_Ixcw4_regx1x : DFFR_X1 port map( D => CU_Ixcw3_1_port, CK => Clk, RN => 
                           n1743, Q => WB_MUX_SEL_MEM_i, QN => n1334);
   CU_Ixcw3_regx6x : DFFR_X1 port map( D => CU_Ixcw2_6_port, CK => Clk, RN => 
                           n1744, Q => PC_SEL_i, QN => n_1106);
   CU_Ixcw2_i_regx11x : DFFR_X1 port map( D => CU_Ixcw1_6_port, CK => Clk, RN 
                           => n1744, Q => CU_Ixcw2_i_11_port, QN => n_1107);
   CU_Ixcw2_i_regx10x : DFFR_X1 port map( D => CU_Ixcw1_10_port, CK => Clk, RN 
                           => n1744, Q => CU_Ixcw2_i_10_port, QN => n_1108);
   DATAPATH_IxSecond_stxIMM_out_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_4_port, CK => Clk,
                           Q => n_1109, QN => n1192);
   DATAPATH_IxSecond_stxIMM_out_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_3_port, CK => Clk,
                           Q => n_1110, QN => n1196);
   DATAPATH_IxSecond_stxIMM_out_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_2_port, CK => Clk,
                           Q => n_1111, QN => n1195);
   DATAPATH_IxSecond_stxIMM_out_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_1_port, CK => Clk,
                           Q => n_1112, QN => n1194);
   DATAPATH_IxSecond_stxIMM_out_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_31_port, CK => Clk
                           , Q => n_1113, QN => n1170);
   DATAPATH_IxSecond_stxIMM_out_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_30_port, CK => Clk
                           , Q => n_1114, QN => n1169);
   DATAPATH_IxSecond_stxIMM_out_regx29x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_29_port, CK => Clk
                           , Q => n_1115, QN => n1157);
   DATAPATH_IxSecond_stxIMM_out_regx28x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_28_port, CK => Clk
                           , Q => n_1116, QN => n1166);
   DATAPATH_IxSecond_stxIMM_out_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_27_port, CK => Clk
                           , Q => n_1117, QN => n1167);
   DATAPATH_IxSecond_stxIMM_out_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_26_port, CK => Clk
                           , Q => n_1118, QN => n1168);
   DATAPATH_IxSecond_stxIMM_out_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_25_port, CK => Clk
                           , Q => n_1119, QN => n1171);
   DATAPATH_IxSecond_stxIMM_out_regx24x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_24_port, CK => Clk
                           , Q => n_1120, QN => n1172);
   DATAPATH_IxSecond_stxIMM_out_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_23_port, CK => Clk
                           , Q => n_1121, QN => n1174);
   DATAPATH_IxSecond_stxIMM_out_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_22_port, CK => Clk
                           , Q => n_1122, QN => n1179);
   DATAPATH_IxSecond_stxIMM_out_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_21_port, CK => Clk
                           , Q => n_1123, QN => n1173);
   DATAPATH_IxSecond_stxIMM_out_regx20x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_20_port, CK => Clk
                           , Q => n_1124, QN => n1178);
   DATAPATH_IxSecond_stxIMM_out_regx19x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_19_port, CK => Clk
                           , Q => n_1125, QN => n1177);
   DATAPATH_IxSecond_stxIMM_out_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_18_port, CK => Clk
                           , Q => n_1126, QN => n1175);
   DATAPATH_IxSecond_stxIMM_out_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_17_port, CK => Clk
                           , Q => n_1127, QN => n1176);
   DATAPATH_IxSecond_stxIMM_out_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_16_port, CK => Clk
                           , Q => n_1128, QN => n1180);
   DATAPATH_IxSecond_stxIMM_out_regx15x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_15_port, CK => Clk
                           , Q => n_1129, QN => n1181);
   DATAPATH_IxSecond_stxIMM_out_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_14_port, CK => Clk
                           , Q => n_1130, QN => n1183);
   DATAPATH_IxSecond_stxIMM_out_regx13x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_13_port, CK => Clk
                           , Q => n_1131, QN => n1188);
   DATAPATH_IxSecond_stxIMM_out_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_12_port, CK => Clk
                           , Q => n_1132, QN => n1182);
   DATAPATH_IxSecond_stxIMM_out_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_0_port, CK => Clk,
                           Q => n_1133, QN => n1193);
   CU_Ixcw3_regx0x : DFFR_X1 port map( D => CU_Ixcw2_0_port, CK => Clk, RN => 
                           n1744, Q => CU_Ixcw3_0_port, QN => n_1134);
   CU_Ixcw4_regx0x : DFFR_X1 port map( D => CU_Ixcw3_0_port, CK => Clk, RN => 
                           n1744, Q => RF_WE_MEM_i, QN => n1333);
   CU_Ixcw5_regx0x : DFFR_X1 port map( D => RF_WE_MEM_i, CK => Clk, RN => n1744
                           , Q => RF_WR_EN, QN => n1299);
   DATAPATH_IxFirst_stxPC_regx1x : DFF_X1 port map( D => n1546, CK => Clk, Q =>
                           DATAPATH_IxPC4_1_port, QN => n1388);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx1x : DFF_X1 port map( D => n1513, CK =>
                           Clk, Q => n1612, QN => n1339);
   DATAPATH_IxSecond_stxPC_out_regx1x : DFF_X1 port map( D => n1512, CK => Clk,
                           Q => n_1135, QN => n1599);
   DATAPATH_IxSecond_stxBR_target_regx1x : DFF_X1 port map( D => n1845, CK => 
                           Clk, Q => n_1136, QN => n1214);
   DATAPATH_IxFirst_stxPC_regx0x : DFF_X1 port map( D => n1547, CK => Clk, Q =>
                           DATAPATH_IxPC4_0_port, QN => n1387);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx0x : DFF_X1 port map( D => n1515, CK =>
                           Clk, Q => DATAPATH_IxSecond_stxjump_target_0_port, 
                           QN => n1338);
   DATAPATH_IxSecond_stxBR_target_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_0_port, CK => Clk, 
                           Q => n_1137, QN => n1213);
   DATAPATH_IxSecond_stxPC_out_regx0x : DFF_X1 port map( D => n1514, CK => Clk,
                           Q => n_1138, QN => n1598);
   DATAPATH_IxFirst_stxPC_regx2x : DFF_X1 port map( D => n1545, CK => Clk, Q =>
                           IRAM_ADD_2_port, QN => n1389);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx2x : DFF_X1 port map( D => n1511, CK =>
                           Clk, Q => n1241, QN => n1610);
   DATAPATH_IxSecond_stxPC_out_regx2x : DFF_X1 port map( D => n1510, CK => Clk,
                           Q => n_1139, QN => n1579);
   DATAPATH_IxSecond_stxBR_target_regx2x : DFF_X1 port map( D => n1296, CK => 
                           Clk, Q => DATAPATH_IxSecond_stxBR_target_2_port, QN 
                           => n_1140);
   DATAPATH_IxFirst_stxPC_regx3x : DFF_X1 port map( D => n1544, CK => Clk, Q =>
                           IRAM_ADD_3_port, QN => n1390);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx3x : DFF_X1 port map( D => n1509, CK =>
                           Clk, Q => n1614, QN => n1340);
   DATAPATH_IxSecond_stxPC_out_regx3x : DFF_X1 port map( D => n1508, CK => Clk,
                           Q => n_1141, QN => n1597);
   DATAPATH_IxSecond_stxBR_target_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_3_port, CK => Clk, 
                           Q => n_1142, QN => n1215);
   DATAPATH_IxFirst_stxPC_regx4x : DFF_X1 port map( D => n1543, CK => Clk, Q =>
                           IRAM_ADD_4_port, QN => n1391);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx4x : DFF_X1 port map( D => n1507, CK =>
                           Clk, Q => n1244, QN => n1620);
   DATAPATH_IxSecond_stxPC_out_regx4x : DFF_X1 port map( D => n1506, CK => Clk,
                           Q => n_1143, QN => n1581);
   DATAPATH_IxSecond_stxBR_target_regx4x : DFF_X1 port map( D => n1839, CK => 
                           Clk, Q => n_1144, QN => n1216);
   DATAPATH_IxFirst_stxPC_regx5x : DFF_X1 port map( D => n1542, CK => Clk, Q =>
                           IRAM_ADD_5_port, QN => n1392);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx5x : DFF_X1 port map( D => n1505, CK =>
                           Clk, Q => n_1145, QN => n1341);
   DATAPATH_IxSecond_stxBR_target_regx5x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_5_port, CK => Clk, 
                           Q => n_1146, QN => n1217);
   DATAPATH_IxSecond_stxPC_out_regx5x : DFF_X1 port map( D => n1504, CK => Clk,
                           Q => n_1147, QN => n1596);
   DATAPATH_IxFirst_stxPC_regx6x : DFF_X1 port map( D => n1541, CK => Clk, Q =>
                           IRAM_ADD_6_port, QN => n1393);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx6x : DFF_X1 port map( D => n1503, CK =>
                           Clk, Q => n_1148, QN => n1342);
   DATAPATH_IxSecond_stxBR_target_regx6x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_6_port, CK => Clk, 
                           Q => DATAPATH_IxSecond_stxBR_target_6_port, QN => 
                           n_1149);
   DATAPATH_IxSecond_stxPC_out_regx6x : DFF_X1 port map( D => n1502, CK => Clk,
                           Q => n_1150, QN => n1595);
   DATAPATH_IxFirst_stxPC_regx7x : DFF_X1 port map( D => n1540, CK => Clk, Q =>
                           IRAM_ADD_7_port, QN => n1394);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx7x : DFF_X1 port map( D => n1501, CK =>
                           Clk, Q => n1248, QN => n1611);
   DATAPATH_IxSecond_stxBR_target_regx7x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_7_port, CK => Clk, 
                           Q => n_1151, QN => n1218);
   DATAPATH_IxSecond_stxPC_out_regx7x : DFF_X1 port map( D => n1500, CK => Clk,
                           Q => n_1152, QN => n1578);
   DATAPATH_IxFirst_stxPC_regx8x : DFF_X1 port map( D => n1539, CK => Clk, Q =>
                           IRAM_ADD_8_port, QN => n1395);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx8x : DFF_X1 port map( D => n1499, CK =>
                           Clk, Q => n_1153, QN => n1343);
   DATAPATH_IxSecond_stxPC_out_regx8x : DFF_X1 port map( D => n1498, CK => Clk,
                           Q => n_1154, QN => n1592);
   DATAPATH_IxSecond_stxBR_target_regx8x : DFF_X1 port map( D => n1291, CK => 
                           Clk, Q => DATAPATH_IxSecond_stxBR_target_8_port, QN 
                           => n_1155);
   DATAPATH_IxFirst_stxPC_regx9x : DFF_X1 port map( D => n1538, CK => Clk, Q =>
                           IRAM_ADD_9_port, QN => n1396);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx9x : DFF_X1 port map( D => n1497, CK =>
                           Clk, Q => n_1156, QN => n1344);
   DATAPATH_IxSecond_stxPC_out_regx9x : DFF_X1 port map( D => n1496, CK => Clk,
                           Q => n_1157, QN => n1594);
   DATAPATH_IxSecond_stxBR_target_regx9x : DFF_X1 port map( D => n1836, CK => 
                           Clk, Q => n_1158, QN => n1219);
   DATAPATH_IxFirst_stxPC_regx10x : DFF_X1 port map( D => n1537, CK => Clk, Q 
                           => IRAM_ADD_10_port, QN => n1397);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx10x : DFF_X1 port map( D => n1495, CK 
                           => Clk, Q => n_1159, QN => n1345);
   DATAPATH_IxSecond_stxPC_out_regx10x : DFF_X1 port map( D => n1494, CK => Clk
                           , Q => n_1160, QN => n1607);
   DATAPATH_IxSecond_stxBR_target_regx10x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_10_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_10_port, QN => 
                           n_1161);
   DATAPATH_IxFirst_stxPC_regx11x : DFF_X1 port map( D => n1536, CK => Clk, Q 
                           => IRAM_ADD_11_port, QN => n1398);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx11x : DFF_X1 port map( D => n1493, CK 
                           => Clk, Q => n_1162, QN => n1346);
   DATAPATH_IxSecond_stxBR_target_regx11x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_11_port, CK => Clk,
                           Q => n_1163, QN => n1220);
   DATAPATH_IxSecond_stxPC_out_regx11x : DFF_X1 port map( D => n1492, CK => Clk
                           , Q => n_1164, QN => n1601);
   DATAPATH_IxFirst_stxPC_regx12x : DFF_X1 port map( D => n1535, CK => Clk, Q 
                           => IRAM_ADD_12_port, QN => n1399);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx12x : DFF_X1 port map( D => n1491, CK 
                           => Clk, Q => n_1165, QN => n1347);
   DATAPATH_IxSecond_stxPC_out_regx12x : DFF_X1 port map( D => n1490, CK => Clk
                           , Q => n_1166, QN => n1606);
   DATAPATH_IxSecond_stxBR_target_regx13x : DFF_X1 port map( D => n1822, CK => 
                           Clk, Q => n_1167, QN => n1221);
   DATAPATH_IxFirst_stxPC_regx13x : DFF_X1 port map( D => n1534, CK => Clk, Q 
                           => IRAM_ADD_13_port, QN => n1400);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx13x : DFF_X1 port map( D => n1489, CK 
                           => Clk, Q => n_1168, QN => n1348);
   DATAPATH_IxSecond_stxPC_out_regx13x : DFF_X1 port map( D => n1488, CK => Clk
                           , Q => n_1169, QN => n1605);
   DATAPATH_IxFirst_stxPC_regx14x : DFF_X1 port map( D => n1533, CK => Clk, Q 
                           => IRAM_ADD_14_port, QN => n1401);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx14x : DFF_X1 port map( D => n1487, CK 
                           => Clk, Q => n1622, QN => n1349);
   DATAPATH_IxSecond_stxPC_out_regx14x : DFF_X1 port map( D => n1486, CK => Clk
                           , Q => n_1170, QN => n1602);
   DATAPATH_IxSecond_stxBR_target_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_14_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_14_port, QN => 
                           n_1171);
   DATAPATH_IxFirst_stxPC_regx15x : DFF_X1 port map( D => n1532, CK => Clk, Q 
                           => IRAM_ADD_15_port, QN => n1402);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx15x : DFF_X1 port map( D => n1485, CK 
                           => Clk, Q => n1257, QN => n1616);
   DATAPATH_IxSecond_stxPC_out_regx15x : DFF_X1 port map( D => n1484, CK => Clk
                           , Q => n_1172, QN => n1580);
   DATAPATH_IxSecond_stxBR_target_regx15x : DFF_X1 port map( D => n1820, CK => 
                           Clk, Q => n_1173, QN => n1222);
   DATAPATH_IxSecond_stxBR_target_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_12_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_12_port, QN => 
                           n_1174);
   DATAPATH_IxSecond_stxBR_target_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_16_port, CK => Clk,
                           Q => n_1175, QN => n1223);
   DATAPATH_IxFirst_stxPC_regx16x : DFF_X1 port map( D => n1531, CK => Clk, Q 
                           => IRAM_ADD_16_port, QN => n1403);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx16x : DFF_X1 port map( D => n1483, CK 
                           => Clk, Q => n_1176, QN => n1350);
   DATAPATH_IxSecond_stxPC_out_regx16x : DFF_X1 port map( D => n1482, CK => Clk
                           , Q => n_1177, QN => n1593);
   DATAPATH_IxSecond_stxBR_target_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_17_port, CK => Clk,
                           Q => n_1178, QN => n1224);
   DATAPATH_IxFirst_stxPC_regx17x : DFF_X1 port map( D => n1530, CK => Clk, Q 
                           => IRAM_ADD_17_port, QN => n1404);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx17x : DFF_X1 port map( D => n1481, CK 
                           => Clk, Q => n_1179, QN => n1351);
   DATAPATH_IxSecond_stxPC_out_regx17x : DFF_X1 port map( D => n1480, CK => Clk
                           , Q => n_1180, QN => n1604);
   DATAPATH_IxSecond_stxBR_target_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_18_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_18_port, QN => 
                           n_1181);
   DATAPATH_IxFirst_stxPC_regx18x : DFF_X1 port map( D => n1529, CK => Clk, Q 
                           => IRAM_ADD_18_port, QN => n1405);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx18x : DFF_X1 port map( D => n1479, CK 
                           => Clk, Q => n_1182, QN => n1352);
   DATAPATH_IxSecond_stxPC_out_regx18x : DFF_X1 port map( D => n1478, CK => Clk
                           , Q => n_1183, QN => n1603);
   DATAPATH_IxFirst_stxPC_regx19x : DFF_X1 port map( D => n1528, CK => Clk, Q 
                           => IRAM_ADD_19_port, QN => n1406);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx19x : DFF_X1 port map( D => n1477, CK 
                           => Clk, Q => n_1184, QN => n1353);
   DATAPATH_IxSecond_stxBR_target_regx19x : DFF_X1 port map( D => n1802, CK => 
                           Clk, Q => n_1185, QN => n1225);
   DATAPATH_IxSecond_stxPC_out_regx19x : DFF_X1 port map( D => n1476, CK => Clk
                           , Q => n_1186, QN => n1600);
   DATAPATH_IxFirst_stxPC_regx20x : DFF_X1 port map( D => n1527, CK => Clk, Q 
                           => IRAM_ADD_20_port, QN => n1407);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx20x : DFF_X1 port map( D => n1475, CK 
                           => Clk, Q => n_1187, QN => n1354);
   DATAPATH_IxSecond_stxPC_out_regx20x : DFF_X1 port map( D => n1474, CK => Clk
                           , Q => n_1188, QN => n1577);
   DATAPATH_IxSecond_stxBR_target_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_21_port, CK => Clk,
                           Q => n_1189, QN => n1227);
   DATAPATH_IxFirst_stxPC_regx21x : DFF_X1 port map( D => n1526, CK => Clk, Q 
                           => IRAM_ADD_21_port, QN => n1408);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx21x : DFF_X1 port map( D => n1473, CK 
                           => Clk, Q => n_1190, QN => n1355);
   DATAPATH_IxSecond_stxPC_out_regx21x : DFF_X1 port map( D => n1472, CK => Clk
                           , Q => n_1191, QN => n1583);
   DATAPATH_IxSecond_stxBR_target_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_22_port, CK => Clk,
                           Q => n_1192, QN => n1228);
   DATAPATH_IxFirst_stxPC_regx22x : DFF_X1 port map( D => n1525, CK => Clk, Q 
                           => IRAM_ADD_22_port, QN => n1409);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx22x : DFF_X1 port map( D => n1471, CK 
                           => Clk, Q => n1619, QN => n1356);
   DATAPATH_IxSecond_stxPC_out_regx22x : DFF_X1 port map( D => n1470, CK => Clk
                           , Q => n_1193, QN => n1586);
   DATAPATH_IxSecond_stxBR_target_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_23_port, CK => Clk,
                           Q => n_1194, QN => n1229);
   DATAPATH_IxFirst_stxPC_regx23x : DFF_X1 port map( D => n1524, CK => Clk, Q 
                           => IRAM_ADD_23_port, QN => n1410);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx23x : DFF_X1 port map( D => n1469, CK 
                           => Clk, Q => n_1195, QN => n1357);
   DATAPATH_IxSecond_stxPC_out_regx23x : DFF_X1 port map( D => n1468, CK => Clk
                           , Q => n_1196, QN => n1588);
   DATAPATH_IxSecond_stxBR_target_regx20x : DFF_X1 port map( D => n1292, CK => 
                           Clk, Q => n_1197, QN => n1226);
   DATAPATH_IxSecond_stxBR_target_regx24x : DFF_X1 port map( D => n1806, CK => 
                           Clk, Q => n_1198, QN => n1230);
   DATAPATH_IxFirst_stxPC_regx24x : DFF_X1 port map( D => n1523, CK => Clk, Q 
                           => IRAM_ADD_24_port, QN => n1411);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx24x : DFF_X1 port map( D => n1467, CK 
                           => Clk, Q => n_1199, QN => n1358);
   DATAPATH_IxSecond_stxPC_out_regx24x : DFF_X1 port map( D => n1466, CK => Clk
                           , Q => n_1200, QN => n1576);
   DATAPATH_IxSecond_stxBR_target_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_25_port, CK => Clk,
                           Q => n_1201, QN => n1231);
   DATAPATH_IxFirst_stxPC_regx25x : DFF_X1 port map( D => n1522, CK => Clk, Q 
                           => IRAM_ADD_25_port, QN => n1412);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx25x : DFF_X1 port map( D => n1465, CK 
                           => Clk, Q => n_1202, QN => n1359);
   DATAPATH_IxSecond_stxPC_out_regx25x : DFF_X1 port map( D => n1464, CK => Clk
                           , Q => n_1203, QN => n1582);
   DATAPATH_IxFirst_stxPC_regx26x : DFF_X1 port map( D => n1521, CK => Clk, Q 
                           => IRAM_ADD_26_port, QN => n1413);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx26x : DFF_X1 port map( D => n1463, CK 
                           => Clk, Q => n1618, QN => n1360);
   DATAPATH_IxSecond_stxPC_out_regx26x : DFF_X1 port map( D => n1462, CK => Clk
                           , Q => n_1204, QN => n1585);
   DATAPATH_IxSecond_stxBR_target_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_26_port, CK => Clk,
                           Q => n_1205, QN => n1232);
   DATAPATH_IxFirst_stxPC_regx27x : DFF_X1 port map( D => n1520, CK => Clk, Q 
                           => IRAM_ADD_27_port, QN => n1414);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx27x : DFF_X1 port map( D => n1461, CK 
                           => Clk, Q => n_1206, QN => n1361);
   DATAPATH_IxSecond_stxBR_target_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_27_port, CK => Clk,
                           Q => n_1207, QN => n1233);
   DATAPATH_IxSecond_stxPC_out_regx27x : DFF_X1 port map( D => n1460, CK => Clk
                           , Q => n_1208, QN => n1587);
   DATAPATH_IxFirst_stxPC_regx28x : DFF_X1 port map( D => n1519, CK => Clk, Q 
                           => IRAM_ADD_28_port, QN => n1415);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx28x : DFF_X1 port map( D => n1459, CK 
                           => Clk, Q => n_1209, QN => n1362);
   DATAPATH_IxSecond_stxPC_out_regx28x : DFF_X1 port map( D => n1458, CK => Clk
                           , Q => n_1210, QN => n1575);
   DATAPATH_IxSecond_stxBR_target_regx29x : DFF_X1 port map( D => n1814, CK => 
                           Clk, Q => n_1211, QN => n1235);
   DATAPATH_IxFirst_stxPC_regx29x : DFF_X1 port map( D => n1518, CK => Clk, Q 
                           => IRAM_ADD_29_port, QN => n1416);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx29x : DFF_X1 port map( D => n1457, CK 
                           => Clk, Q => n_1212, QN => n1363);
   DATAPATH_IxSecond_stxPC_out_regx29x : DFF_X1 port map( D => n1456, CK => Clk
                           , Q => n_1213, QN => n1574);
   DATAPATH_IxSecond_stxBR_target_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_30_port, CK => Clk,
                           Q => n_1214, QN => n1236);
   DATAPATH_IxFirst_stxPC_regx30x : DFF_X1 port map( D => n1517, CK => Clk, Q 
                           => IRAM_ADD_30_port, QN => n1417);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx30x : DFF_X1 port map( D => n1455, CK 
                           => Clk, Q => n1617, QN => n1364);
   DATAPATH_IxSecond_stxPC_out_regx30x : DFF_X1 port map( D => n1454, CK => Clk
                           , Q => n_1215, QN => n1584);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_1_port, CK => Clk, Q 
                           => DRAM_ADD_1_port, QN => n1420);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx1x : DFF_X1 port map( D => 
                           DRAM_ADD_1_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_1_port, QN => n_1216);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_2_port, CK => Clk, Q 
                           => DRAM_ADD_2_port, QN => n1421);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx2x : DFF_X1 port map( D => 
                           DRAM_ADD_2_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_2_port, QN => n_1217);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_3_port, CK => Clk, Q 
                           => DRAM_ADD_3_port, QN => n1422);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx3x : DFF_X1 port map( D => 
                           DRAM_ADD_3_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_3_port, QN => n_1218);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_4_port, CK => Clk, Q 
                           => DRAM_ADD_4_port, QN => n1423);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx4x : DFF_X1 port map( D => 
                           DRAM_ADD_4_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_4_port, QN => n_1219);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx5x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_5_port, CK => Clk, Q 
                           => DRAM_ADD_5_port, QN => n1424);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx5x : DFF_X1 port map( D => 
                           DRAM_ADD_5_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_5_port, QN => n_1220);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx6x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_6_port, CK => Clk, Q 
                           => DRAM_ADD_6_port, QN => n1425);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx6x : DFF_X1 port map( D => 
                           DRAM_ADD_6_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_6_port, QN => n_1221);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx7x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_7_port, CK => Clk, Q 
                           => DRAM_ADD_7_port, QN => n1426);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx7x : DFF_X1 port map( D => 
                           DRAM_ADD_7_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_7_port, QN => n_1222);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx8x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_8_port, CK => Clk, Q 
                           => DRAM_ADD_8_port, QN => n1427);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx8x : DFF_X1 port map( D => 
                           DRAM_ADD_8_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_8_port, QN => n_1223);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx9x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_9_port, CK => Clk, Q 
                           => DRAM_ADD_9_port, QN => n1428);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx9x : DFF_X1 port map( D => 
                           DRAM_ADD_9_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_9_port, QN => n_1224);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx11x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_11_port, CK => Clk, Q 
                           => DRAM_ADD_11_port, QN => n1430);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx11x : DFF_X1 port map( D => 
                           DRAM_ADD_11_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_11_port, QN => n_1225);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_12_port, CK => Clk, Q 
                           => DRAM_ADD_12_port, QN => n1431);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx12x : DFF_X1 port map( D => 
                           DRAM_ADD_12_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_12_port, QN => n_1226);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx13x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_13_port, CK => Clk, Q 
                           => DRAM_ADD_13_port, QN => n1432);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx13x : DFF_X1 port map( D => 
                           DRAM_ADD_13_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_13_port, QN => n_1227);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_14_port, CK => Clk, Q 
                           => DRAM_ADD_14_port, QN => n1433);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx14x : DFF_X1 port map( D => 
                           DRAM_ADD_14_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_14_port, QN => n_1228);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx15x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_15_port, CK => Clk, Q 
                           => DRAM_ADD_15_port, QN => n1434);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx15x : DFF_X1 port map( D => 
                           DRAM_ADD_15_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_15_port, QN => n_1229);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx19x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_19_port, CK => Clk, Q 
                           => DRAM_ADD_19_port, QN => n1438);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx19x : DFF_X1 port map( D => 
                           DRAM_ADD_19_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_19_port, QN => n_1230);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx20x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_20_port, CK => Clk, Q 
                           => DRAM_ADD_20_port, QN => n1439);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx20x : DFF_X1 port map( D => 
                           DRAM_ADD_20_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_20_port, QN => n_1231);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_21_port, CK => Clk, Q 
                           => DRAM_ADD_21_port, QN => n1440);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx21x : DFF_X1 port map( D => 
                           DRAM_ADD_21_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_21_port, QN => n_1232);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_22_port, CK => Clk, Q 
                           => DRAM_ADD_22_port, QN => n1441);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx22x : DFF_X1 port map( D => 
                           DRAM_ADD_22_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_22_port, QN => n_1233);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_23_port, CK => Clk, Q 
                           => DRAM_ADD_23_port, QN => n1442);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx23x : DFF_X1 port map( D => 
                           DRAM_ADD_23_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_23_port, QN => n_1234);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx24x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_24_port, CK => Clk, Q 
                           => DRAM_ADD_24_port, QN => n1443);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx24x : DFF_X1 port map( D => 
                           DRAM_ADD_24_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_24_port, QN => n_1235);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_27_port, CK => Clk, Q 
                           => DRAM_ADD_27_port, QN => n1446);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx27x : DFF_X1 port map( D => 
                           DRAM_ADD_27_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_27_port, QN => n_1236);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx28x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_28_port, CK => Clk, Q 
                           => DRAM_ADD_28_port, QN => n1447);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx28x : DFF_X1 port map( D => 
                           DRAM_ADD_28_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_28_port, QN => n_1237);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx29x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_29_port, CK => Clk, Q 
                           => DRAM_ADD_29_port, QN => n1448);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx29x : DFF_X1 port map( D => 
                           DRAM_ADD_29_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_29_port, QN => n_1238);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_30_port, CK => Clk, Q 
                           => DRAM_ADD_30_port, QN => n1449);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx30x : DFF_X1 port map( D => 
                           DRAM_ADD_30_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_30_port, QN => n_1239);
   DATAPATH_IxSecond_stxBR_target_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_31_port, CK => Clk,
                           Q => n_1240, QN => n1237);
   DATAPATH_IxFirst_stxPC_regx31x : DFF_X1 port map( D => n1516, CK => Clk, Q 
                           => IRAM_ADD_31_port, QN => n1418);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx31x : DFF_X1 port map( D => n1453, CK 
                           => Clk, Q => n_1241, QN => n1365);
   DATAPATH_IxSecond_stxPC_out_regx31x : DFF_X1 port map( D => n1452, CK => Clk
                           , Q => n_1242, QN => n1589);
   DATAPATH_IxSecond_stxBR_target_regx28x : DFF_X1 port map( D => n1811, CK => 
                           Clk, Q => n_1243, QN => n1234);
   U5 : NAND3_X1 port map( A1 => n22, A2 => n23, A3 => n1754, ZN => n1287);
   U10 : NAND3_X1 port map( A1 => n32, A2 => n33, A3 => n1755, ZN => n1288);
   U13 : NAND3_X1 port map( A1 => n33, A2 => n23, A3 => n36, ZN => n1289);
   U19 : NAND3_X1 port map( A1 => IRAM_DOUT(14), A2 => IRAM_DOUT(12), A3 => n43
                           , ZN => n32);
   U22 : NAND3_X1 port map( A1 => IRAM_DOUT(5), A2 => n28, A3 => IRAM_DOUT(2), 
                           ZN => n33);
   U115 : NAND3_X1 port map( A1 => IRAM_ADD_28_port, A2 => IRAM_ADD_27_port, A3
                           => n118, ZN => n110);
   U124 : XOR2_X1 port map( A => n1815, B => n126, Z => n47);
   U153 : XOR2_X1 port map( A => n1810, B => n152, Z => n46);
   U165 : XOR2_X1 port map( A => n1409, B => n164, Z => n162);
   U182 : XOR2_X1 port map( A => n180, B => n181, Z => n1292);
   U280 : XOR2_X1 port map( A => n268, B => n269, Z => n48);
   U304 : NAND3_X1 port map( A1 => n1852, A2 => n165, A3 => n1744, ZN => n289);
   U387 : XOR2_X1 port map( A => n358, B => n359, Z => n356);
   U389 : XOR2_X1 port map( A => n363, B => n359, Z => n355);
   U397 : XOR2_X1 port map( A => n360, B => n375, Z => n374);
   U399 : XOR2_X1 port map( A => n364, B => n375, Z => n373);
   U404 : XOR2_X1 port map( A => n386, B => n387, Z => n383);
   U416 : XOR2_X1 port map( A => n403, B => n404, Z => n402);
   U430 : XOR2_X1 port map( A => n432, B => n433, Z => n431);
   U431 : XOR2_X1 port map( A => n434, B => n433, Z => n428);
   U457 : XOR2_X1 port map( A => n474, B => n475, Z => n473);
   U459 : XOR2_X1 port map( A => n479, B => n475, Z => n470);
   U467 : XOR2_X1 port map( A => n476, B => n491, Z => n490);
   U469 : NAND3_X1 port map( A1 => n1863, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, A3 => n495, ZN 
                           => n493);
   U471 : XOR2_X1 port map( A => n480, B => n491, Z => n489);
   U477 : XOR2_X1 port map( A => n504, B => n505, Z => n501);
   U491 : XOR2_X1 port map( A => n523, B => n524, Z => n522);
   U493 : XOR2_X1 port map( A => n528, B => n524, Z => n519);
   U500 : XOR2_X1 port map( A => n525, B => n539, Z => n538);
   U502 : NAND3_X1 port map( A1 => n1867, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, A3 => n543, ZN 
                           => n541);
   U504 : XOR2_X1 port map( A => n529, B => n539, Z => n537);
   U510 : XOR2_X1 port map( A => n552, B => n553, Z => n549);
   U523 : XOR2_X1 port map( A => n442, B => n568, Z => n567);
   U533 : XOR2_X1 port map( A => n581, B => n582, Z => n579);
   U535 : XOR2_X1 port map( A => n586, B => n582, Z => n578);
   U542 : XOR2_X1 port map( A => n583, B => n597, Z => n596);
   U545 : XOR2_X1 port map( A => n587, B => n597, Z => n595);
   U566 : XOR2_X1 port map( A => n629, B => n630, Z => n628);
   U568 : XOR2_X1 port map( A => n634, B => n630, Z => n625);
   U575 : XOR2_X1 port map( A => n631, B => n645, Z => n644);
   U577 : XOR2_X1 port map( A => n635, B => n645, Z => n643);
   U582 : XOR2_X1 port map( A => n656, B => n657, Z => n653);
   U594 : XOR2_X1 port map( A => n673, B => n674, Z => n672);
   U596 : XOR2_X1 port map( A => n678, B => n674, Z => n671);
   U603 : XOR2_X1 port map( A => n675, B => n689, Z => n688);
   U606 : XOR2_X1 port map( A => n679, B => n689, Z => n687);
   U608 : NAND3_X1 port map( A1 => n1880, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, A3 => n337, ZN 
                           => n693);
   U615 : NAND3_X1 port map( A1 => n1335, A2 => n1673, A3 => n1336, ZN => n418)
                           ;
   U625 : XOR2_X1 port map( A => n420, B => n707, Z => n706);
   U626 : XOR2_X1 port map( A => n708, B => n709, Z => n707);
   U628 : XOR2_X1 port map( A => n420, B => n712, Z => n710);
   U629 : XOR2_X1 port map( A => n708, B => n713, Z => n712);
   U695 : XOR2_X1 port map( A => n1664, B => n655, Z => n657);
   U699 : XOR2_X1 port map( A => n1664, B => n1916, Z => n658);
   U710 : XOR2_X1 port map( A => n1664, B => n333, Z => n336);
   U725 : XOR2_X1 port map( A => n1664, B => n1734, Z => n388);
   U727 : XOR2_X1 port map( A => n1664, B => n399, Z => n404);
   U740 : XOR2_X1 port map( A => n1664, B => n438, Z => n441);
   U750 : XOR2_X1 port map( A => n1664, B => n663, Z => n664);
   U767 : XOR2_X1 port map( A => n1664, B => n610, Z => n783);
   U783 : XOR2_X1 port map( A => n791, B => n792, Z => n237);
   U787 : XOR2_X1 port map( A => n798, B => n799, Z => n797);
   U789 : XOR2_X1 port map( A => n803, B => n799, Z => n795);
   U794 : XOR2_X1 port map( A => n800, B => n808, Z => n807);
   U796 : XOR2_X1 port map( A => n804, B => n808, Z => n806);
   U798 : XOR2_X1 port map( A => n812, B => n813, Z => 
                           DATAPATH_IxSecond_stxjump_target_5_port);
   U804 : XOR2_X1 port map( A => n821, B => n822, Z => n820);
   U806 : XOR2_X1 port map( A => n825, B => n822, Z => n818);
   U807 : XOR2_X1 port map( A => n1365, B => n1386, Z => n822);
   U811 : XOR2_X1 port map( A => n829, B => n824, Z => n828);
   U813 : XOR2_X1 port map( A => n826, B => n829, Z => n827);
   U834 : XOR2_X1 port map( A => n838, B => n843, Z => n847);
   U836 : XOR2_X1 port map( A => n845, B => n838, Z => n846);
   U856 : XOR2_X1 port map( A => n854, B => n860, Z => n864);
   U858 : XOR2_X1 port map( A => n862, B => n854, Z => n863);
   U872 : XOR2_X1 port map( A => n879, B => n869, Z => n182);
   U888 : XOR2_X1 port map( A => n898, B => n874, Z => 
                           DATAPATH_IxSecond_stxjump_target_17_port);
   U915 : XOR2_X1 port map( A => n905, B => n910, Z => n920);
   U917 : XOR2_X1 port map( A => n905, B => n917, Z => n918);
   U937 : XOR2_X1 port map( A => n1384, B => n1343, Z => n244);
   U946 : XOR2_X1 port map( A => n940, B => n930, Z => n939);
   U948 : XOR2_X1 port map( A => n944, B => n930, Z => n938);
   U955 : XOR2_X1 port map( A => n942, B => n931, Z => n948);
   U958 : XOR2_X1 port map( A => n946, B => n931, Z => n947);
   U963 : NAND3_X1 port map( A1 => n1343, A2 => n1962, A3 => n1384, ZN => n951)
                           ;
   U969 : XOR2_X1 port map( A => n1383, B => n1248, Z => n799);
   U985 : XOR2_X1 port map( A => n958, B => n1340, Z => n815);
   U999 : XOR2_X1 port map( A => n1382, B => n1342, Z => n808);
   U1192 : XOR2_X1 port map( A => n1897, B => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, Z => n463);
   U1296 : XOR2_X1 port map( A => n1741, B => 
                           DATAPATH_IxThird_stxALU_IN1_0_port, Z => n700);
   U1341 : NAND3_X1 port map( A1 => n1673, A2 => n1591, A3 => n1335, ZN => n790
                           );
   U1353 : XOR2_X1 port map( A => n1739, B => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, Z => n565);
   U1368 : XOR2_X1 port map( A => n1149, B => n1165, Z => n1097);
   U1370 : XOR2_X1 port map( A => n1151, B => n1161, Z => n1101);
   U1371 : XOR2_X1 port map( A => n1148, B => n1162, Z => n1100);
   U1372 : XOR2_X1 port map( A => n1147, B => n1163, Z => n1099);
   U1373 : XOR2_X1 port map( A => n1150, B => n1164, Z => n1098);
   U1376 : XOR2_X1 port map( A => n1158, B => n1164, Z => n1107);
   U1377 : XOR2_X1 port map( A => n1160, B => n1165, Z => n1106);
   U1398 : XOR2_X1 port map( A => n1149, B => n1156, Z => n1121);
   U1400 : XOR2_X1 port map( A => n1151, B => n1152, Z => n1125);
   U1401 : XOR2_X1 port map( A => n1147, B => n1153, Z => n1124);
   U1402 : XOR2_X1 port map( A => n1150, B => n1154, Z => n1123);
   U1403 : XOR2_X1 port map( A => n1148, B => n1155, Z => n1122);
   U1407 : XOR2_X1 port map( A => n1155, B => n1159, Z => n1131);
   U1408 : XOR2_X1 port map( A => n1156, B => n1160, Z => n1130);
   U1422 : NAND3_X1 port map( A1 => n1134, A2 => n26, A3 => n1139, ZN => 
                           CU_IxN24);
   U310 : NOR3_X2 port map( A1 => n1745, A2 => n109, A3 => n165, ZN => n190);
   DATAPATH_IxSecond_stxIMM_out_regx11x : DFF_X1 port map( D => n1631, CK => 
                           Clk, Q => n_1244, QN => n1187);
   DATAPATH_IxSecond_stxIMM_out_regx10x : DFF_X1 port map( D => n1630, CK => 
                           Clk, Q => n_1245, QN => n1186);
   DATAPATH_IxSecond_stxIMM_out_regx9x : DFF_X1 port map( D => n1629, CK => Clk
                           , Q => n_1246, QN => n1184);
   DATAPATH_IxSecond_stxIMM_out_regx8x : DFF_X1 port map( D => n1628, CK => Clk
                           , Q => n_1247, QN => n1185);
   DATAPATH_IxSecond_stxIMM_out_regx7x : DFF_X1 port map( D => n1627, CK => Clk
                           , Q => n_1248, QN => n1189);
   DATAPATH_IxSecond_stxIMM_out_regx6x : DFF_X1 port map( D => n1626, CK => Clk
                           , Q => n_1249, QN => n1190);
   DATAPATH_IxSecond_stxIMM_out_regx5x : DFF_X1 port map( D => n1625, CK => Clk
                           , Q => n_1250, QN => n1191);
   CU_Ixcw5_regx1x : DFFR_X1 port map( D => WB_MUX_SEL_MEM_i, CK => Clk, RN => 
                           n1744, Q => n1682, QN => n1573);
   CU_Ixstate_var_regx0x : DFFR_X1 port map( D => CU_IxN51, CK => Clk, RN => 
                           n1743, Q => n_1251, QN => n1298);
   CU_Ixstate_var_regx1x : DFFR_X1 port map( D => CU_IxN52, CK => Clk, RN => 
                           n1744, Q => n1923, QN => n1197);
   CU_Ixcw2_i_regx14x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1743, Q => n_1252, QN => n1211);
   CU_Ixcw2_i_regx13x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1743, Q => n_1253, QN => n1212);
   CU_Ixcw2_i_regx8x : DFFR_X1 port map( D => CU_Ixcw1_8_port, CK => Clk, RN =>
                           n1743, Q => n_1254, QN => n1206);
   CU_Ixcw2_i_regx7x : DFFR_X1 port map( D => CU_Ixcw1_7_port, CK => Clk, RN =>
                           n1744, Q => n_1255, QN => n1207);
   CU_Ixcw2_i_regx5x : DFFR_X1 port map( D => CU_Ixcw1_5_port, CK => Clk, RN =>
                           n1744, Q => n_1256, QN => n1203);
   CU_Ixcw2_i_regx4x : DFFR_X1 port map( D => CU_Ixcw1_4_port, CK => Clk, RN =>
                           n1744, Q => n_1257, QN => n1202);
   CU_Ixcw2_i_regx2x : DFFR_X1 port map( D => CU_Ixcw1_2_port, CK => Clk, RN =>
                           n1744, Q => n_1258, QN => n1200);
   CU_Ixcw2_i_regx1x : DFFR_X1 port map( D => CU_Ixcw1_1_port, CK => Clk, RN =>
                           n1744, Q => n_1259, QN => n1199);
   CU_Ixcw2_i_regx0x : DFFR_X1 port map( D => CU_Ixcw1_0_port, CK => Clk, RN =>
                           n1744, Q => n_1260, QN => n1198);
   CU_Ixcw2_i_regx9x : DFFR_X1 port map( D => CU_Ixcw1_9_port, CK => Clk, RN =>
                           n1744, Q => n_1261, QN => n1205);
   CU_Ixcw2_i_regx6x : DFFR_X1 port map( D => CU_Ixcw1_6_port, CK => Clk, RN =>
                           n1744, Q => n_1262, QN => n1204);
   CU_Ixcw2_i_regx3x : DFFR_X1 port map( D => CU_Ixcw1_9_port, CK => Clk, RN =>
                           n1744, Q => n_1263, QN => n1201);
   U1445 : INV_X1 port map( A => n1113, ZN => n1966);
   U1446 : INV_X1 port map( A => n1090, ZN => n1968);
   U1447 : OAI221_X1 port map( B1 => n1703, B2 => n1574, C1 => n1448, C2 => 
                           n1700, A => n1032, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_29_port);
   U1448 : OAI221_X1 port map( B1 => n1703, B2 => n1575, C1 => n1447, C2 => 
                           n1700, A => n1029, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_28_port);
   U1449 : OAI221_X1 port map( B1 => n1702, B2 => n1576, C1 => n1443, C2 => 
                           n1699, A => n1019, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_24_port);
   U1450 : OAI221_X1 port map( B1 => n1702, B2 => n1577, C1 => n1439, C2 => 
                           n1699, A => n994, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_20_port);
   U1451 : OAI221_X1 port map( B1 => n1703, B2 => n1592, C1 => n1427, C2 => 
                           n1700, A => n1037, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_8_port);
   U1452 : NOR3_X1 port map( A1 => n1746, A2 => n109, A3 => n1852, ZN => n191);
   U1453 : AOI211_X2 port map( C1 => n1923, C2 => n1298, A => n1747, B => n296,
                           ZN => n109);
   U1454 : OAI221_X1 port map( B1 => n1702, B2 => n1593, C1 => n1435, C2 => 
                           n1699, A => n991, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_16_port);
   U1455 : OR2_X1 port map( A1 => n1636, A2 => n1335, ZN => n1590);
   U1456 : NOR2_X1 port map( A1 => n1849, A2 => n1381, ZN => n1625);
   U1457 : NOR2_X1 port map( A1 => n1849, A2 => n1382, ZN => n1626);
   U1458 : NOR2_X1 port map( A1 => n1849, A2 => n1383, ZN => n1627);
   U1459 : NOR2_X1 port map( A1 => n1849, A2 => n1384, ZN => n1628);
   U1460 : NOR2_X1 port map( A1 => n1849, A2 => n1624, ZN => n1629);
   U1461 : NOR2_X1 port map( A1 => n1849, A2 => n1385, ZN => n1630);
   U1462 : NOR2_X1 port map( A1 => n1386, A2 => n1849, ZN => n1631);
   U1463 : OR4_X1 port map( A1 => n1746, A2 => n109, A3 => n159, A4 => n1851, 
                           ZN => n108);
   U1464 : INV_X1 port map( A => n108, ZN => n1632);
   U1465 : NOR3_X1 port map( A1 => n1854, A2 => n1211, A3 => n291, ZN => n159);
   U1466 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_1_port, Z => n1739
                           );
   U1467 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_0_port, Z => n1741
                           );
   U1468 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_3_port, Z => n1735
                           );
   U1469 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_2_port, Z => n1737
                           );
   U1470 : INV_X1 port map( A => n441, ZN => n1888);
   U1471 : NOR2_X1 port map( A1 => n1655, A2 => n1664, ZN => n401);
   U1472 : INV_X1 port map( A => n571, ZN => n1926);
   U1473 : INV_X1 port map( A => n882, ZN => n1830);
   U1474 : OAI22_X1 port map( A1 => n1860, A2 => n725, B1 => n726, B2 => n429, 
                           ZN => n420);
   U1475 : XNOR2_X1 port map( A => n709, B => n717, ZN => n726);
   U1476 : XNOR2_X1 port map( A => n713, B => n717, ZN => n725);
   U1477 : BUF_X1 port map( A => n979, Z => n1694);
   U1478 : BUF_X1 port map( A => n985, Z => n1683);
   U1479 : BUF_X1 port map( A => n985, Z => n1684);
   U1480 : BUF_X1 port map( A => n979, Z => n1695);
   U1481 : BUF_X1 port map( A => n985, Z => n1685);
   U1482 : BUF_X1 port map( A => n979, Z => n1696);
   U1483 : INV_X1 port map( A => n429, ZN => n1860);
   U1484 : INV_X1 port map( A => n1673, ZN => n1663);
   U1485 : INV_X1 port map( A => n1672, ZN => n1662);
   U1486 : INV_X1 port map( A => n1673, ZN => n1664);
   U1487 : BUF_X1 port map( A => n108, Z => n1646);
   U1488 : BUF_X1 port map( A => n108, Z => n1644);
   U1489 : BUF_X1 port map( A => n108, Z => n1645);
   U1490 : BUF_X1 port map( A => n1766, Z => n1649);
   U1491 : BUF_X1 port map( A => n1766, Z => n1650);
   U1492 : INV_X1 port map( A => n783, ZN => n1871);
   U1493 : XNOR2_X1 port map( A => n1667, B => n422, ZN => n717);
   U1494 : XNOR2_X1 port map( A => n1337, B => n1856, ZN => n454);
   U1495 : AOI21_X1 port map( B1 => n364, B2 => n361, A => n362, ZN => n363);
   U1496 : BUF_X1 port map( A => n299, Z => n1713);
   U1497 : AOI21_X1 port map( B1 => n635, B2 => n632, A => n633, ZN => n634);
   U1498 : BUF_X1 port map( A => n1765, Z => n1648);
   U1499 : AOI21_X1 port map( B1 => n360, B2 => n361, A => n362, ZN => n358);
   U1500 : BUF_X1 port map( A => n54, Z => n1717);
   U1501 : BUF_X1 port map( A => n54, Z => n1718);
   U1502 : BUF_X1 port map( A => n1765, Z => n1647);
   U1503 : BUF_X1 port map( A => n299, Z => n1712);
   U1504 : BUF_X1 port map( A => n54, Z => n1719);
   U1505 : AOI21_X1 port map( B1 => n412, B2 => n406, A => n407, ZN => n411);
   U1506 : AOI22_X1 port map( A1 => n1886, A2 => n373, B1 => n374, B2 => n357, 
                           ZN => n367);
   U1507 : XNOR2_X1 port map( A => n405, B => n441, ZN => n440);
   U1508 : AOI21_X1 port map( B1 => n587, B2 => n584, A => n585, ZN => n586);
   U1509 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n633, ZN => n629);
   U1510 : AOI21_X1 port map( B1 => n405, B2 => n406, A => n407, ZN => n403);
   U1511 : INV_X1 port map( A => n357, ZN => n1886);
   U1512 : INV_X1 port map( A => n464, ZN => n1859);
   U1513 : BUF_X1 port map( A => n1928, Z => n1654);
   U1514 : BUF_X1 port map( A => n1928, Z => n1655);
   U1515 : NOR2_X1 port map( A1 => n1672, A2 => n1655, ZN => n571);
   U1516 : BUF_X1 port map( A => n1928, Z => n1656);
   U1517 : OAI22_X1 port map( A1 => n1861, A2 => n737, B1 => n738, B2 => n475, 
                           ZN => n429);
   U1518 : XNOR2_X1 port map( A => n1662, B => n1898, ZN => n737);
   U1519 : AOI21_X1 port map( B1 => n491, B2 => n739, A => n478, ZN => n738);
   U1520 : OAI21_X1 port map( B1 => n740, B2 => n505, A => n492, ZN => n739);
   U1521 : OAI22_X1 port map( A1 => n1887, A2 => n778, B1 => n779, B2 => n404, 
                           ZN => n357);
   U1522 : XNOR2_X1 port map( A => n1665, B => n1735, ZN => n778);
   U1523 : AOI21_X1 port map( B1 => n1888, B2 => n780, A => n407, ZN => n779);
   U1524 : OAI21_X1 port map( B1 => n781, B2 => n568, A => n444, ZN => n780);
   U1525 : NOR2_X1 port map( A1 => n1847, A2 => n882, ZN => n896);
   U1526 : INV_X1 port map( A => n1681, ZN => n1674);
   U1527 : NOR2_X1 port map( A1 => n1847, A2 => n1386, ZN => n882);
   U1528 : XNOR2_X1 port map( A => n1666, B => n565, ZN => n568);
   U1529 : XNOR2_X1 port map( A => n1893, B => DATAPATH_IxThird_stxALU1xN222, 
                           ZN => n422);
   U1530 : XNOR2_X1 port map( A => n1662, B => n700, ZN => n696);
   U1531 : XNOR2_X1 port map( A => n1737, B => n1889, ZN => n438);
   U1532 : OAI22_X1 port map( A1 => n1819, A2 => n889, B1 => n876, B2 => n890, 
                           ZN => DATAPATH_IxSecond_stxjump_target_18_port);
   U1533 : XNOR2_X1 port map( A => n870, B => n886, ZN => n889);
   U1534 : XNOR2_X1 port map( A => n870, B => n885, ZN => n890);
   U1535 : XNOR2_X1 port map( A => n1735, B => n1887, ZN => n399);
   U1536 : NOR2_X1 port map( A1 => n413, A2 => n1889, ZN => n407);
   U1537 : BUF_X1 port map( A => n975, Z => n1702);
   U1538 : BUF_X1 port map( A => n975, Z => n1703);
   U1539 : INV_X1 port map( A => n1634, ZN => n1687);
   U1540 : INV_X1 port map( A => n1634, ZN => n1686);
   U1541 : INV_X1 port map( A => n1633, ZN => n1698);
   U1542 : INV_X1 port map( A => n1633, ZN => n1697);
   U1543 : XNOR2_X1 port map( A => n1663, B => n393, ZN => n394);
   U1544 : BUF_X1 port map( A => n982, Z => n1688);
   U1545 : BUF_X1 port map( A => n982, Z => n1689);
   U1546 : BUF_X1 port map( A => n976, Z => n1699);
   U1547 : BUF_X1 port map( A => n976, Z => n1700);
   U1548 : BUF_X1 port map( A => n981, Z => n1691);
   U1549 : BUF_X1 port map( A => n981, Z => n1692);
   U1550 : XNOR2_X1 port map( A => n1663, B => n1739, ZN => n447);
   U1551 : XNOR2_X1 port map( A => n1663, B => n1741, ZN => n569);
   U1552 : XNOR2_X1 port map( A => n1663, B => n1730, ZN => n380);
   U1553 : BUF_X1 port map( A => n976, Z => n1701);
   U1554 : XNOR2_X1 port map( A => n1666, B => n1737, ZN => n413);
   U1555 : BUF_X1 port map( A => n981, Z => n1693);
   U1556 : INV_X1 port map( A => n626, ZN => n1877);
   U1557 : NAND4_X1 port map( A1 => n1871, A2 => n580, A3 => n597, A4 => n755, 
                           ZN => n754);
   U1558 : NOR2_X1 port map( A1 => n582, A2 => n619, ZN => n755);
   U1559 : BUF_X1 port map( A => n975, Z => n1704);
   U1560 : AOI21_X1 port map( B1 => n696, B2 => n1671, A => n1892, ZN => n781);
   U1561 : INV_X1 port map( A => n446, ZN => n1892);
   U1562 : BUF_X1 port map( A => n982, Z => n1690);
   U1563 : OAI21_X1 port map( B1 => n1876, B2 => n657, A => n648, ZN => n759);
   U1564 : INV_X1 port map( A => n763, ZN => n1876);
   U1565 : OAI21_X1 port map( B1 => n664, B2 => n1877, A => n647, ZN => n763);
   U1566 : OAI21_X1 port map( B1 => n776, B2 => n387, A => n378, ZN => n775);
   U1567 : AOI21_X1 port map( B1 => n394, B2 => n357, A => n1885, ZN => n776);
   U1568 : INV_X1 port map( A => n379, ZN => n1885);
   U1569 : NOR2_X1 port map( A1 => n469, A2 => n487, ZN => n1022);
   U1570 : AND3_X1 port map( A1 => n1701, A2 => n1633, A3 => n1704, ZN => n979)
                           ;
   U1571 : AND3_X1 port map( A1 => n1634, A2 => n1690, A3 => n1693, ZN => n985)
                           ;
   U1572 : OR4_X1 port map( A1 => n512, A2 => n503, A3 => n422, A4 => n427, ZN 
                           => n972);
   U1573 : INV_X1 port map( A => n876, ZN => n1819);
   U1574 : OR4_X1 port map( A1 => n353, A2 => n655, A3 => n669, A4 => n686, ZN 
                           => n1035);
   U1575 : INV_X1 port map( A => n452, ZN => n1856);
   U1576 : NAND2_X1 port map( A1 => n1819, A2 => n1825, ZN => n900);
   U1577 : OR3_X1 port map( A1 => n663, A2 => n624, A3 => n642, ZN => n1036);
   U1578 : INV_X1 port map( A => n182, ZN => n1802);
   U1579 : INV_X1 port map( A => n46, ZN => n1806);
   U1580 : INV_X1 port map( A => n1728, ZN => n1720);
   U1581 : XNOR2_X1 port map( A => n1662, B => n594, ZN => n597);
   U1582 : XNOR2_X1 port map( A => n1665, B => n576, ZN => n582);
   U1583 : XNOR2_X1 port map( A => n1670, B => n624, ZN => n630);
   U1584 : XNOR2_X1 port map( A => n1670, B => n669, ZN => n674);
   U1585 : XNOR2_X1 port map( A => n1671, B => n353, ZN => n359);
   U1586 : NOR2_X1 port map( A1 => n365, A2 => n1884, ZN => n362);
   U1587 : NOR2_X1 port map( A1 => n588, A2 => n1870, ZN => n585);
   U1588 : NOR2_X1 port map( A1 => n680, A2 => n1879, ZN => n677);
   U1589 : NOR2_X1 port map( A1 => n636, A2 => n1875, ZN => n633);
   U1590 : XNOR2_X1 port map( A => n1664, B => n642, ZN => n645);
   U1591 : XNOR2_X1 port map( A => n1664, B => n686, ZN => n689);
   U1592 : XNOR2_X1 port map( A => n1664, B => n371, ZN => n375);
   U1593 : XNOR2_X1 port map( A => n1669, B => n618, ZN => n619);
   U1594 : XNOR2_X1 port map( A => n1664, B => n347, ZN => n348);
   U1595 : XNOR2_X1 port map( A => n1662, B => n560, ZN => n561);
   U1596 : AOI22_X1 port map( A1 => n613, A2 => n1872, B1 => n1912, B2 => n1873
                           , ZN => n611);
   U1597 : NAND2_X1 port map( A1 => n601, A2 => n580, ZN => n613);
   U1598 : XNOR2_X1 port map( A => n1666, B => n385, ZN => n387);
   U1599 : AOI22_X1 port map( A1 => n489, A2 => n471, B1 => n1864, B2 => n490, 
                           ZN => n483);
   U1600 : INV_X1 port map( A => n190, ZN => n1766);
   U1601 : INV_X1 port map( A => n520, ZN => n1868);
   U1602 : INV_X1 port map( A => n580, ZN => n1873);
   U1603 : INV_X1 port map( A => n471, ZN => n1864);
   U1604 : AOI21_X1 port map( B1 => n647, B2 => n1877, A => n649, ZN => n656);
   U1605 : BUF_X1 port map( A => n1613, Z => n1673);
   U1606 : NOR2_X1 port map( A1 => n1971, A2 => n1645, ZN => n168);
   U1607 : BUF_X1 port map( A => n1669, Z => n1672);
   U1608 : BUF_X1 port map( A => n1670, Z => n1667);
   U1609 : BUF_X1 port map( A => n1670, Z => n1665);
   U1610 : BUF_X1 port map( A => n1668, Z => n1666);
   U1611 : BUF_X1 port map( A => n1670, Z => n1671);
   U1612 : INV_X1 port map( A => n48, ZN => n1839);
   U1613 : INV_X1 port map( A => n49, ZN => n1845);
   U1614 : INV_X1 port map( A => n206, ZN => n1820);
   U1615 : INV_X1 port map( A => n217, ZN => n1822);
   U1616 : XNOR2_X1 port map( A => n1668, B => n518, ZN => n524);
   U1617 : NOR2_X1 port map( A1 => n481, A2 => n1862, ZN => n478);
   U1618 : XNOR2_X1 port map( A => n1667, B => n469, ZN => n475);
   U1619 : NOR2_X1 port map( A1 => n530, A2 => n1866, ZN => n527);
   U1620 : XNOR2_X1 port map( A => n1337, B => n427, ZN => n433);
   U1621 : XNOR2_X1 port map( A => n1662, B => n536, ZN => n539);
   U1622 : XNOR2_X1 port map( A => n1662, B => n487, ZN => n491);
   U1623 : XNOR2_X1 port map( A => n1337, B => n463, ZN => n464);
   U1624 : AOI21_X1 port map( B1 => n679, B2 => n676, A => n677, ZN => n678);
   U1625 : XNOR2_X1 port map( A => n1662, B => n512, ZN => n513);
   U1626 : AOI21_X1 port map( B1 => n476, B2 => n477, A => n478, ZN => n474);
   U1627 : AOI21_X1 port map( B1 => n525, B2 => n526, A => n527, ZN => n523);
   U1628 : AOI21_X1 port map( B1 => n434, B2 => n727, A => n719, ZN => n713);
   U1629 : AOI21_X1 port map( B1 => n432, B2 => n727, A => n719, ZN => n709);
   U1630 : AOI21_X1 port map( B1 => n480, B2 => n477, A => n478, ZN => n479);
   U1631 : AOI21_X1 port map( B1 => n529, B2 => n526, A => n527, ZN => n528);
   U1632 : BUF_X1 port map( A => n92, Z => n1714);
   U1633 : BUF_X1 port map( A => n92, Z => n1715);
   U1634 : BUF_X1 port map( A => n1757, Z => n1642);
   U1635 : BUF_X1 port map( A => n1757, Z => n1641);
   U1636 : BUF_X1 port map( A => n1757, Z => n1643);
   U1637 : OAI21_X1 port map( B1 => n443, B2 => n446, A => n444, ZN => n412);
   U1638 : OAI21_X1 port map( B1 => n442, B2 => n443, A => n444, ZN => n405);
   U1639 : XNOR2_X1 port map( A => n1669, B => n551, ZN => n553);
   U1640 : XNOR2_X1 port map( A => n1668, B => n503, ZN => n505);
   U1641 : OAI21_X1 port map( B1 => n646, B2 => n647, A => n648, ZN => n631);
   U1642 : OAI21_X1 port map( B1 => n377, B2 => n379, A => n378, ZN => n364);
   U1643 : OAI21_X1 port map( B1 => n649, B2 => n646, A => n648, ZN => n635);
   U1644 : OAI21_X1 port map( B1 => n376, B2 => n377, A => n378, ZN => n360);
   U1645 : INV_X1 port map( A => n191, ZN => n1765);
   U1646 : AOI21_X1 port map( B1 => n1886, B2 => n379, A => n376, ZN => n386);
   U1647 : INV_X1 port map( A => n338, ZN => n1882);
   U1648 : AOI21_X1 port map( B1 => n583, B2 => n584, A => n585, ZN => n581);
   U1649 : AOI21_X1 port map( B1 => n675, B2 => n676, A => n677, ZN => n673);
   U1650 : NAND2_X1 port map( A1 => n1743, A2 => n1714, ZN => n299);
   U1651 : NAND2_X1 port map( A1 => n1643, A2 => n1743, ZN => n54);
   U1652 : INV_X1 port map( A => CU_IxN25, ZN => n1751);
   U1653 : OAI211_X1 port map( C1 => n395, C2 => n1926, A => n397, B => n398, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_3_port);
   U1654 : XNOR2_X1 port map( A => n404, B => n411, ZN => n395);
   U1655 : AOI22_X1 port map( A1 => n400, A2 => n1735, B1 => n401, B2 => n402, 
                           ZN => n397);
   U1656 : AOI22_X1 port map( A1 => n1651, A2 => n399, B1 => 
                           DATAPATH_IxThird_stxALU1xN194, B2 => n1711, ZN => 
                           n398);
   U1657 : INV_X1 port map( A => n729, ZN => n1896);
   U1658 : OAI211_X1 port map( C1 => n435, C2 => n1926, A => n436, B => n437, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_2_port);
   U1659 : XNOR2_X1 port map( A => n412, B => n1888, ZN => n435);
   U1660 : AOI22_X1 port map( A1 => n439, A2 => n1737, B1 => n401, B2 => n440, 
                           ZN => n436);
   U1661 : AOI22_X1 port map( A1 => n1651, A2 => n438, B1 => 
                           DATAPATH_IxThird_stxALU1xN193, B2 => n1711, ZN => 
                           n437);
   U1662 : OAI211_X1 port map( C1 => n1926, C2 => n562, A => n563, B => n564, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_1_port);
   U1663 : XNOR2_X1 port map( A => n446, B => n568, ZN => n562);
   U1664 : AOI22_X1 port map( A1 => n1890, A2 => n1739, B1 => n401, B2 => n567,
                           ZN => n563);
   U1665 : AOI22_X1 port map( A1 => n1652, A2 => n565, B1 => 
                           DATAPATH_IxThird_stxALU1xN192, B2 => n1709, ZN => 
                           n564);
   U1666 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU1xN222, Z => n1638);
   U1667 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU1xN222, Z => n1637);
   U1668 : BUF_X1 port map( A => n1637, Z => n1639);
   U1669 : INV_X1 port map( A => n463, ZN => n1858);
   U1670 : NAND2_X1 port map( A1 => n481, A2 => n1862, ZN => n477);
   U1671 : NAND2_X1 port map( A1 => n365, A2 => n1884, ZN => n361);
   U1672 : NAND2_X1 port map( A1 => n413, A2 => n1889, ZN => n406);
   U1673 : NAND2_X1 port map( A1 => n530, A2 => n1866, ZN => n526);
   U1674 : NAND2_X1 port map( A1 => n588, A2 => n1870, ZN => n584);
   U1675 : NAND2_X1 port map( A1 => n636, A2 => n1875, ZN => n632);
   U1676 : NAND2_X1 port map( A1 => n680, A2 => n1879, ZN => n676);
   U1677 : BUF_X1 port map( A => n1613, Z => n1668);
   U1678 : BUF_X1 port map( A => n1613, Z => n1670);
   U1679 : BUF_X1 port map( A => n1613, Z => n1669);
   U1680 : INV_X1 port map( A => n601, ZN => n1912);
   U1681 : INV_X1 port map( A => n732, ZN => n1857);
   U1682 : NAND2_X1 port map( A1 => n600, A2 => n602, ZN => n587);
   U1683 : OR3_X1 port map( A1 => n599, A2 => n1872, A3 => n1912, ZN => n602);
   U1684 : BUF_X1 port map( A => n92, Z => n1716);
   U1685 : AND2_X1 port map( A1 => CU_Ixcw_LUT_6_port, A2 => n1853, ZN => 
                           CU_Ixcw1_6_port);
   U1686 : INV_X1 port map( A => n1749, ZN => CU_Ixcw_LUT_6_port);
   U1687 : AND2_X1 port map( A1 => CU_Ixcw_LUT_9_port, A2 => n1853, ZN => 
                           CU_Ixcw1_9_port);
   U1688 : AND2_X1 port map( A1 => CU_Ixcw_LUT_10_port, A2 => n1853, ZN => 
                           CU_Ixcw1_10_port);
   U1689 : INV_X1 port map( A => n1590, ZN => n1705);
   U1690 : INV_X1 port map( A => n1590, ZN => n1706);
   U1691 : BUF_X1 port map( A => n1925, Z => n1651);
   U1692 : BUF_X1 port map( A => n1925, Z => n1652);
   U1693 : BUF_X1 port map( A => n1925, Z => n1653);
   U1694 : INV_X1 port map( A => n421, ZN => n1928);
   U1695 : INV_X1 port map( A => n28, ZN => n1756);
   U1696 : OAI221_X1 port map( B1 => n751, B2 => n582, C1 => n1869, C2 => n753,
                           A => n754, ZN => n520);
   U1697 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_19_port, ZN => 
                           n1869);
   U1698 : XNOR2_X1 port map( A => n1664, B => n1908, ZN => n753);
   U1699 : AOI21_X1 port map( B1 => n597, B2 => n784, A => n585, ZN => n751);
   U1700 : OAI22_X1 port map( A1 => n1865, A2 => n744, B1 => n745, B2 => n524, 
                           ZN => n471);
   U1701 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_23_port, ZN => 
                           n1865);
   U1702 : XNOR2_X1 port map( A => n1662, B => n1903, ZN => n744);
   U1703 : AOI21_X1 port map( B1 => n539, B2 => n746, A => n527, ZN => n745);
   U1704 : OAI22_X1 port map( A1 => n1874, A2 => n757, B1 => n758, B2 => n630, 
                           ZN => n580);
   U1705 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_15_port, ZN => 
                           n1874);
   U1706 : XNOR2_X1 port map( A => n1664, B => n1913, ZN => n757);
   U1707 : AOI21_X1 port map( B1 => n645, B2 => n759, A => n633, ZN => n758);
   U1708 : OAI22_X1 port map( A1 => n1616, A2 => n1824, B1 => n903, B2 => n904,
                           ZN => n876);
   U1709 : INV_X1 port map( A => n913, ZN => n1824);
   U1710 : AOI21_X1 port map( B1 => n905, B2 => n906, A => n907, ZN => n903);
   U1711 : OAI21_X1 port map( B1 => n1831, B2 => n909, A => n910, ZN => n906);
   U1712 : OAI22_X1 port map( A1 => n1878, A2 => n765, B1 => n766, B2 => n674, 
                           ZN => n626);
   U1713 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_11_port, ZN => 
                           n1878);
   U1714 : XNOR2_X1 port map( A => n1664, B => n1917, ZN => n765);
   U1715 : AOI21_X1 port map( B1 => n689, B2 => n767, A => n677, ZN => n766);
   U1716 : NAND2_X1 port map( A1 => n1827, A2 => n884, ZN => n879);
   U1717 : OAI211_X1 port map( C1 => n885, C2 => n876, A => n886, B => n887, ZN
                           => n884);
   U1718 : INV_X1 port map( A => n1732, ZN => n1730);
   U1719 : XNOR2_X1 port map( A => n1920, B => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, ZN => n347);
   U1720 : XNOR2_X1 port map( A => n1734, B => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, ZN => n393);
   U1721 : INV_X1 port map( A => n897, ZN => n1847);
   U1722 : XNOR2_X1 port map( A => n1732, B => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, ZN => n385);
   U1723 : XNOR2_X1 port map( A => n372, B => n1884, ZN => n371);
   U1724 : XNOR2_X1 port map( A => n1914, B => 
                           DATAPATH_IxThird_stxALU_IN1_14_port, ZN => n642);
   U1725 : XNOR2_X1 port map( A => n488, B => n1862, ZN => n487);
   U1726 : XNOR2_X1 port map( A => n1913, B => 
                           DATAPATH_IxThird_stxALU_IN1_15_port, ZN => n624);
   U1727 : XNOR2_X1 port map( A => n789, B => n1861, ZN => n469);
   U1728 : NAND2_X1 port map( A1 => n877, A2 => n900, ZN => n898);
   U1729 : XNOR2_X1 port map( A => n1901, B => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, ZN => n512);
   U1730 : XNOR2_X1 port map( A => n1906, B => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n560);
   U1731 : AOI21_X1 port map( B1 => n911, B2 => n921, A => n922, ZN => n910);
   U1732 : XNOR2_X1 port map( A => n1911, B => 
                           DATAPATH_IxThird_stxALU_IN1_16_port, ZN => n618);
   U1733 : XNOR2_X1 port map( A => n1921, B => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, ZN => n353);
   U1734 : XNOR2_X1 port map( A => n1900, B => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, ZN => n503);
   U1735 : XNOR2_X1 port map( A => n1905, B => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, ZN => n551);
   U1736 : XNOR2_X1 port map( A => n1909, B => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, ZN => n594);
   U1737 : XNOR2_X1 port map( A => n1903, B => 
                           DATAPATH_IxThird_stxALU_IN1_23_port, ZN => n518);
   U1738 : XNOR2_X1 port map( A => n1904, B => 
                           DATAPATH_IxThird_stxALU_IN1_22_port, ZN => n536);
   U1739 : XNOR2_X1 port map( A => n1917, B => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, ZN => n669);
   U1740 : XNOR2_X1 port map( A => n1894, B => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, ZN => n427);
   U1741 : XNOR2_X1 port map( A => n1908, B => 
                           DATAPATH_IxThird_stxALU_IN1_19_port, ZN => n576);
   U1742 : XNOR2_X1 port map( A => n1918, B => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, ZN => n686);
   U1743 : XNOR2_X1 port map( A => n1919, B => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, ZN => n333);
   U1744 : INV_X1 port map( A => n326, ZN => n1853);
   U1745 : XNOR2_X1 port map( A => n1916, B => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, ZN => n663);
   U1746 : OAI22_X1 port map( A1 => n1810, A2 => n840, B1 => n835, B2 => n841, 
                           ZN => DATAPATH_IxSecond_stxjump_target_27_port);
   U1747 : XNOR2_X1 port map( A => n844, B => n839, ZN => n840);
   U1748 : XNOR2_X1 port map( A => n834, B => n839, ZN => n841);
   U1749 : OAI21_X1 port map( B1 => n1660, B2 => n1618, A => n845, ZN => n844);
   U1750 : OAI22_X1 port map( A1 => n1805, A2 => n863, B1 => n864, B2 => n181, 
                           ZN => DATAPATH_IxSecond_stxjump_target_22_port);
   U1751 : OAI22_X1 port map( A1 => n1805, A2 => n857, B1 => n181, B2 => n858, 
                           ZN => DATAPATH_IxSecond_stxjump_target_23_port);
   U1752 : XNOR2_X1 port map( A => n861, B => n855, ZN => n857);
   U1753 : XNOR2_X1 port map( A => n851, B => n855, ZN => n858);
   U1754 : OAI21_X1 port map( B1 => n1660, B2 => n1619, A => n862, ZN => n861);
   U1755 : OAI22_X1 port map( A1 => n1810, A2 => n846, B1 => n847, B2 => n835, 
                           ZN => DATAPATH_IxSecond_stxjump_target_26_port);
   U1756 : OAI22_X1 port map( A1 => n1729, A2 => n715, B1 => n716, B2 => n717, 
                           ZN => n708);
   U1757 : AOI21_X1 port map( B1 => n433, B2 => n718, A => n719, ZN => n716);
   U1758 : OAI22_X1 port map( A1 => n1855, A2 => n1896, B1 => n722, B2 => n454,
                           ZN => n718);
   U1759 : AOI22_X1 port map( A1 => n1859, A2 => n429, B1 => n457, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, ZN => n722);
   U1760 : XNOR2_X1 port map( A => n1910, B => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, ZN => n610);
   U1761 : XNOR2_X1 port map( A => n1915, B => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n655);
   U1762 : OAI221_X1 port map( B1 => n1893, B2 => n416, C1 => n1801, C2 => n418
                           , A => n419, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_31_port);
   U1763 : AOI21_X1 port map( B1 => n1708, B2 => n1637, A => n1705, ZN => n416)
                           ;
   U1764 : INV_X1 port map( A => n422, ZN => n1801);
   U1765 : AOI22_X1 port map( A1 => n1638, A2 => n1709, B1 => n420, B2 => n421,
                           ZN => n419);
   U1766 : AOI21_X1 port map( B1 => n1610, B2 => n1846, A => n279, ZN => n817);
   U1767 : INV_X1 port map( A => n283, ZN => n1846);
   U1768 : NAND4_X1 port map( A1 => n967, A2 => n968, A3 => n969, A4 => n970, 
                           ZN => n294);
   U1769 : NOR4_X1 port map( A1 => n565, A2 => n399, A3 => n790, A4 => n438, ZN
                           => n967);
   U1770 : NOR4_X1 port map( A1 => n1035, A2 => n1036, A3 => n333, A4 => n347, 
                           ZN => n969);
   U1771 : NOR4_X1 port map( A1 => n371, A2 => n385, A3 => n393, A4 => n700, ZN
                           => n968);
   U1772 : XNOR2_X1 port map( A => n1895, B => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, ZN => n452);
   U1773 : NOR2_X1 port map( A1 => n916, A2 => n907, ZN => n905);
   U1774 : AOI21_X1 port map( B1 => n710, B2 => n429, A => n1591, ZN => n702);
   U1775 : AOI22_X1 port map( A1 => n513, A2 => n471, B1 => n495, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, ZN => n740);
   U1776 : OR2_X1 port map( A1 => n1088, A2 => n1968, ZN => n1633);
   U1777 : OR2_X1 port map( A1 => n1111, A2 => n1966, ZN => n1634);
   U1778 : OAI21_X1 port map( B1 => n1829, B2 => n900, A => n901, ZN => 
                           DATAPATH_IxSecond_stxjump_target_16_port);
   U1779 : OAI21_X1 port map( B1 => n878, B2 => n1829, A => n876, ZN => n901);
   U1780 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_2_port, ZN => 
                           n1889);
   U1781 : NAND2_X1 port map( A1 => n388, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, ZN => n379);
   U1782 : OAI22_X1 port map( A1 => n1883, A2 => n773, B1 => n774, B2 => n359, 
                           ZN => n338);
   U1783 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_7_port, ZN => 
                           n1883);
   U1784 : XNOR2_X1 port map( A => n1664, B => n1921, ZN => n773);
   U1785 : AOI21_X1 port map( B1 => n375, B2 => n775, A => n362, ZN => n774);
   U1786 : NAND2_X1 port map( A1 => n569, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_0_port, ZN => n446);
   U1787 : INV_X1 port map( A => n835, ZN => n1810);
   U1788 : NAND2_X1 port map( A1 => n380, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, ZN => n378);
   U1789 : NAND2_X1 port map( A1 => n447, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, ZN => n444);
   U1790 : INV_X1 port map( A => n819, ZN => n1815);
   U1791 : OAI21_X1 port map( B1 => n769, B2 => n336, A => n692, ZN => n767);
   U1792 : AOI22_X1 port map( A1 => n348, A2 => n338, B1 => n337, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, ZN => n769);
   U1793 : OAI21_X1 port map( B1 => n748, B2 => n553, A => n540, ZN => n746);
   U1794 : AOI22_X1 port map( A1 => n561, A2 => n520, B1 => n543, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n748);
   U1795 : INV_X1 port map( A => n291, ZN => n1850);
   U1796 : INV_X1 port map( A => n181, ZN => n1805);
   U1797 : INV_X1 port map( A => n268, ZN => n1844);
   U1798 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_26_port, ZN => 
                           n1862);
   U1799 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_6_port, ZN => 
                           n1884);
   U1800 : OAI211_X1 port map( C1 => n696, C2 => n1927, A => n698, B => n699, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_0_port);
   U1801 : INV_X1 port map( A => n401, ZN => n1927);
   U1802 : AOI222_X1 port map( A1 => DATAPATH_IxThird_stxALU1xN191, A2 => n1711
                           , B1 => n571, B2 => n696, C1 => n1653, C2 => n700, 
                           ZN => n699);
   U1803 : AOI22_X1 port map( A1 => n702, A2 => n703, B1 => n1891, B2 => n1741,
                           ZN => n698);
   U1804 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_3_port, ZN => 
                           n1887);
   U1805 : NAND2_X1 port map( A1 => n286, A2 => n1612, ZN => n279);
   U1806 : BUF_X1 port map( A => n1682, Z => n1675);
   U1807 : BUF_X1 port map( A => n1682, Z => n1676);
   U1808 : BUF_X1 port map( A => n1682, Z => n1677);
   U1809 : BUF_X1 port map( A => n1682, Z => n1680);
   U1810 : BUF_X1 port map( A => n1682, Z => n1678);
   U1811 : BUF_X1 port map( A => n1682, Z => n1679);
   U1812 : INV_X1 port map( A => n919, ZN => n1831);
   U1813 : NAND2_X1 port map( A1 => n1115, A2 => n1116, ZN => n1113);
   U1814 : NAND2_X1 port map( A1 => n1093, A2 => n1092, ZN => n1090);
   U1815 : BUF_X1 port map( A => n1682, Z => n1681);
   U1816 : OR2_X1 port map( A1 => n1113, A2 => n1111, ZN => n982);
   U1817 : OR2_X1 port map( A1 => n1090, A2 => n1088, ZN => n975);
   U1818 : NAND2_X1 port map( A1 => n1111, A2 => n1113, ZN => n981);
   U1819 : NAND2_X1 port map( A1 => n1088, A2 => n1090, ZN => n976);
   U1820 : INV_X1 port map( A => n271, ZN => n1838);
   U1821 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_27_port, ZN => 
                           n1861);
   U1822 : NAND2_X1 port map( A1 => n911, A2 => n912, ZN => n909);
   U1823 : INV_X1 port map( A => n734, ZN => n1895);
   U1824 : INV_X1 port map( A => n742, ZN => n1901);
   U1825 : INV_X1 port map( A => n749, ZN => n1905);
   U1826 : INV_X1 port map( A => n750, ZN => n1906);
   U1827 : INV_X1 port map( A => n762, ZN => n1915);
   U1828 : INV_X1 port map( A => n770, ZN => n1919);
   U1829 : INV_X1 port map( A => n771, ZN => n1920);
   U1830 : INV_X1 port map( A => n741, ZN => n1900);
   U1831 : INV_X1 port map( A => n787, ZN => n1910);
   U1832 : INV_X1 port map( A => n788, ZN => n1911);
   U1833 : INV_X1 port map( A => n731, ZN => n1894);
   U1834 : INV_X1 port map( A => n747, ZN => n1904);
   U1835 : INV_X1 port map( A => n760, ZN => n1914);
   U1836 : INV_X1 port map( A => n785, ZN => n1909);
   U1837 : INV_X1 port map( A => n768, ZN => n1918);
   U1838 : NAND2_X1 port map( A1 => n817, A2 => n284, ZN => n282);
   U1839 : INV_X1 port map( A => n715, ZN => n1893);
   U1840 : INV_X1 port map( A => n735, ZN => n1897);
   U1841 : INV_X1 port map( A => n47, ZN => n1811);
   U1842 : INV_X1 port map( A => n111, ZN => n1814);
   U1843 : XNOR2_X1 port map( A => n1663, B => n771, ZN => n337);
   U1844 : NOR2_X1 port map( A1 => n270, A2 => n271, ZN => n269);
   U1845 : XNOR2_X1 port map( A => n1662, B => n788, ZN => n601);
   U1846 : XNOR2_X1 port map( A => n904, B => n914, ZN => n206);
   U1847 : NOR2_X1 port map( A1 => n915, A2 => n907, ZN => n914);
   U1848 : AOI211_X1 port map( C1 => n1831, C2 => n910, A => n916, B => n917, 
                           ZN => n915);
   U1849 : OAI21_X1 port map( B1 => n270, B2 => n1844, A => n1838, ZN => n812);
   U1850 : AOI21_X1 port map( B1 => n101, B2 => n1632, A => n109, ZN => n103);
   U1851 : AOI21_X1 port map( B1 => n132, B2 => n1632, A => n109, ZN => n139);
   U1852 : AOI21_X1 port map( B1 => n144, B2 => n1632, A => n109, ZN => n150);
   U1853 : AOI21_X1 port map( B1 => n172, B2 => n1632, A => n109, ZN => n179);
   U1854 : AOI21_X1 port map( B1 => n198, B2 => n1632, A => n109, ZN => n205);
   U1855 : OAI22_X1 port map( A1 => n1831, A2 => n918, B1 => n919, B2 => n920, 
                           ZN => DATAPATH_IxSecond_stxjump_target_14_port);
   U1856 : OAI22_X1 port map( A1 => n1837, A2 => n947, B1 => n948, B2 => n936, 
                           ZN => DATAPATH_IxSecond_stxjump_target_10_port);
   U1857 : OAI22_X1 port map( A1 => n1844, A2 => n806, B1 => n268, B2 => n807, 
                           ZN => DATAPATH_IxSecond_stxjump_target_6_port);
   U1858 : OAI22_X1 port map( A1 => n1837, A2 => n938, B1 => n939, B2 => n936, 
                           ZN => DATAPATH_IxSecond_stxjump_target_11_port);
   U1859 : OAI21_X1 port map( B1 => n941, B2 => n942, A => n1961, ZN => n940);
   U1860 : OAI22_X1 port map( A1 => n795, A2 => n1844, B1 => n268, B2 => n797, 
                           ZN => DATAPATH_IxSecond_stxjump_target_7_port);
   U1861 : OAI21_X1 port map( B1 => n804, B2 => n801, A => n1964, ZN => n803);
   U1862 : INV_X1 port map( A => n1451, ZN => n1849);
   U1863 : OAI221_X1 port map( B1 => n1654, B2 => n514, C1 => n1903, C2 => n516
                           , A => n517, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_23_port);
   U1864 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_23_port, A => n1706, ZN 
                           => n516);
   U1865 : AOI22_X1 port map( A1 => n1652, A2 => n518, B1 => 
                           DATAPATH_IxThird_stxALU1xN214, B2 => n1710, ZN => 
                           n517);
   U1866 : AOI22_X1 port map( A1 => n519, A2 => n520, B1 => n1868, B2 => n522, 
                           ZN => n514);
   U1867 : OAI221_X1 port map( B1 => n1654, B2 => n532, C1 => n1904, C2 => n534
                           , A => n535, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_22_port);
   U1868 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_22_port, A => n1706, ZN 
                           => n534);
   U1869 : AOI22_X1 port map( A1 => n1652, A2 => n536, B1 => 
                           DATAPATH_IxThird_stxALU1xN213, B2 => n1710, ZN => 
                           n535);
   U1870 : AOI22_X1 port map( A1 => n537, A2 => n520, B1 => n1868, B2 => n538, 
                           ZN => n532);
   U1871 : OAI221_X1 port map( B1 => n1654, B2 => n465, C1 => n1898, C2 => n467
                           , A => n468, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_27_port);
   U1872 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_27_port, A => n1705, ZN 
                           => n467);
   U1873 : AOI22_X1 port map( A1 => n1651, A2 => n469, B1 => 
                           DATAPATH_IxThird_stxALU1xN218, B2 => n1710, ZN => 
                           n468);
   U1874 : AOI22_X1 port map( A1 => n470, A2 => n471, B1 => n1864, B2 => n473, 
                           ZN => n465);
   U1875 : OAI221_X1 port map( B1 => n1654, B2 => n483, C1 => n1899, C2 => n485
                           , A => n486, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_26_port);
   U1876 : INV_X1 port map( A => n488, ZN => n1899);
   U1877 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_26_port, A => n1705, ZN 
                           => n485);
   U1878 : AOI22_X1 port map( A1 => n1652, A2 => n487, B1 => 
                           DATAPATH_IxThird_stxALU1xN217, B2 => n1710, ZN => 
                           n486);
   U1879 : OAI221_X1 port map( B1 => n1895, B2 => n449, C1 => n1655, C2 => n450
                           , A => n451, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_29_port);
   U1880 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, A => n1705, ZN 
                           => n449);
   U1881 : AOI22_X1 port map( A1 => n1651, A2 => n452, B1 => 
                           DATAPATH_IxThird_stxALU1xN220, B2 => n1710, ZN => 
                           n451);
   U1882 : XNOR2_X1 port map( A => n453, B => n454, ZN => n450);
   U1883 : OAI221_X1 port map( B1 => n1897, B2 => n459, C1 => n1655, C2 => n460
                           , A => n461, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_28_port);
   U1884 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, A => n1705, ZN 
                           => n459);
   U1885 : AOI22_X1 port map( A1 => n1651, A2 => n1858, B1 => 
                           DATAPATH_IxThird_stxALU1xN219, B2 => n1710, ZN => 
                           n461);
   U1886 : XNOR2_X1 port map( A => n1860, B => n464, ZN => n460);
   U1887 : OAI221_X1 port map( B1 => n1905, B2 => n548, C1 => n1655, C2 => n549
                           , A => n550, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_21_port);
   U1888 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, A => n1706, ZN 
                           => n548);
   U1889 : AOI22_X1 port map( A1 => n1652, A2 => n551, B1 => 
                           DATAPATH_IxThird_stxALU1xN212, B2 => n1710, ZN => 
                           n550);
   U1890 : OAI221_X1 port map( B1 => n1900, B2 => n500, C1 => n1655, C2 => n501
                           , A => n502, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_25_port);
   U1891 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, A => n1706, ZN 
                           => n500);
   U1892 : AOI22_X1 port map( A1 => n1652, A2 => n503, B1 => 
                           DATAPATH_IxThird_stxALU1xN216, B2 => n1710, ZN => 
                           n502);
   U1893 : OAI221_X1 port map( B1 => n1911, B2 => n615, C1 => n1656, C2 => n616
                           , A => n617, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_16_port);
   U1894 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_16_port, A => n1706, ZN 
                           => n615);
   U1895 : AOI22_X1 port map( A1 => n1652, A2 => n618, B1 => 
                           DATAPATH_IxThird_stxALU1xN207, B2 => n1709, ZN => 
                           n617);
   U1896 : XNOR2_X1 port map( A => n1873, B => n619, ZN => n616);
   U1897 : OAI21_X1 port map( B1 => n1829, B2 => n1828, A => n1826, ZN => n886)
                           ;
   U1898 : OAI21_X1 port map( B1 => n1828, B2 => n1825, A => n1826, ZN => n885)
                           ;
   U1899 : OAI221_X1 port map( B1 => n1915, B2 => n652, C1 => n1655, C2 => n653
                           , A => n654, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_13_port);
   U1900 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, A => n1705, ZN 
                           => n652);
   U1901 : AOI22_X1 port map( A1 => n1653, A2 => n655, B1 => 
                           DATAPATH_IxThird_stxALU1xN204, B2 => n1709, ZN => 
                           n654);
   U1902 : INV_X1 port map( A => n965, ZN => n1848);
   U1903 : AOI21_X1 port map( B1 => n962, B2 => n961, A => n1386, ZN => n965);
   U1904 : AOI21_X1 port map( B1 => n912, B2 => n911, A => n922, ZN => n917);
   U1905 : NOR3_X1 port map( A1 => IRAM_ADD_25_port, A2 => n132, A3 => n1644, 
                           ZN => n143);
   U1906 : NOR3_X1 port map( A1 => IRAM_ADD_23_port, A2 => n144, A3 => n1645, 
                           ZN => n156);
   U1907 : XNOR2_X1 port map( A => n1667, B => n372, ZN => n365);
   U1908 : AOI21_X1 port map( B1 => n809, B2 => n1838, A => n811, ZN => n800);
   U1909 : AOI21_X1 port map( B1 => n809, B2 => n270, A => n811, ZN => n804);
   U1910 : XNOR2_X1 port map( A => n1663, B => n770, ZN => n695);
   U1911 : XNOR2_X1 port map( A => n1664, B => n787, ZN => n605);
   U1912 : XNOR2_X1 port map( A => n1663, B => n762, ZN => n650);
   U1913 : XNOR2_X1 port map( A => n1665, B => n785, ZN => n588);
   U1914 : XNOR2_X1 port map( A => n1671, B => n768, ZN => n680);
   U1915 : XNOR2_X1 port map( A => n1670, B => n760, ZN => n636);
   U1916 : XNOR2_X1 port map( A => n924, B => n925, ZN => n217);
   U1917 : NAND2_X1 port map( A1 => n911, A2 => n1823, ZN => n924);
   U1918 : OAI21_X1 port map( B1 => n919, B2 => n921, A => n912, ZN => n925);
   U1919 : INV_X1 port map( A => n922, ZN => n1823);
   U1920 : OAI21_X1 port map( B1 => n286, B2 => n1612, A => n279, ZN => n49);
   U1921 : OAI21_X1 port map( B1 => n118, B2 => n1646, A => n1767, ZN => n124);
   U1922 : OAI21_X1 port map( B1 => n192, B2 => n1646, A => n1767, ZN => n194);
   U1923 : OAI21_X1 port map( B1 => n214, B2 => n1646, A => n1767, ZN => n216);
   U1924 : OAI21_X1 port map( B1 => n224, B2 => n1645, A => n1767, ZN => n226);
   U1925 : OAI21_X1 port map( B1 => n234, B2 => n1646, A => n1767, ZN => n236);
   U1926 : OAI21_X1 port map( B1 => n246, B2 => n1645, A => n1767, ZN => n248);
   U1927 : OAI21_X1 port map( B1 => n256, B2 => n1646, A => n1767, ZN => n258);
   U1928 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_2_port, A => n1767, 
                           ZN => n267);
   U1929 : OAI22_X1 port map( A1 => n1723, A2 => n1578, B1 => n1611, B2 => 
                           n1721, ZN => n1500);
   U1930 : OAI22_X1 port map( A1 => n1722, A2 => n1581, B1 => n1620, B2 => 
                           n1721, ZN => n1506);
   U1931 : OAI22_X1 port map( A1 => n1722, A2 => n1579, B1 => n1610, B2 => 
                           n1721, ZN => n1510);
   U1932 : OAI22_X1 port map( A1 => n1725, A2 => n1580, B1 => n1616, B2 => 
                           n1720, ZN => n1484);
   U1933 : OAI221_X1 port map( B1 => n1654, B2 => n423, C1 => n1894, C2 => n425
                           , A => n426, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_30_port);
   U1934 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, A => n1705, ZN 
                           => n425);
   U1935 : AOI22_X1 port map( A1 => n1651, A2 => n427, B1 => 
                           DATAPATH_IxThird_stxALU1xN221, B2 => n1710, ZN => 
                           n426);
   U1936 : AOI22_X1 port map( A1 => n428, A2 => n429, B1 => n1860, B2 => n431, 
                           ZN => n423);
   U1937 : OAI221_X1 port map( B1 => n1654, B2 => n572, C1 => n1908, C2 => n574
                           , A => n575, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_19_port);
   U1938 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_19_port, A => n1706, ZN 
                           => n574);
   U1939 : AOI22_X1 port map( A1 => n1652, A2 => n576, B1 => 
                           DATAPATH_IxThird_stxALU1xN210, B2 => n1709, ZN => 
                           n575);
   U1940 : AOI22_X1 port map( A1 => n1873, A2 => n578, B1 => n579, B2 => n580, 
                           ZN => n572);
   U1941 : OAI221_X1 port map( B1 => n1654, B2 => n590, C1 => n1909, C2 => n592
                           , A => n593, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_18_port);
   U1942 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, A => n1706, ZN 
                           => n592);
   U1943 : AOI22_X1 port map( A1 => n1652, A2 => n594, B1 => 
                           DATAPATH_IxThird_stxALU1xN209, B2 => n1709, ZN => 
                           n593);
   U1944 : AOI22_X1 port map( A1 => n1873, A2 => n595, B1 => n596, B2 => n580, 
                           ZN => n590);
   U1945 : XNOR2_X1 port map( A => n244, B => n1837, ZN => n1291);
   U1946 : OAI221_X1 port map( B1 => n1906, B2 => n557, C1 => n1655, C2 => n558
                           , A => n559, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_20_port);
   U1947 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, A => n1706, ZN 
                           => n557);
   U1948 : AOI22_X1 port map( A1 => n1652, A2 => n560, B1 => 
                           DATAPATH_IxThird_stxALU1xN211, B2 => n1710, ZN => 
                           n559);
   U1949 : XNOR2_X1 port map( A => n520, B => n561, ZN => n558);
   U1950 : OAI21_X1 port map( B1 => n455, B2 => n429, A => n1857, ZN => n453);
   U1951 : AND2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_28_port, A2 => 
                           n457, ZN => n455);
   U1952 : XNOR2_X1 port map( A => n927, B => n919, ZN => 
                           DATAPATH_IxSecond_stxjump_target_12_port);
   U1953 : NAND2_X1 port map( A1 => n912, A2 => n1821, ZN => n927);
   U1954 : INV_X1 port map( A => n921, ZN => n1821);
   U1955 : INV_X1 port map( A => n936, ZN => n1837);
   U1956 : OAI221_X1 port map( B1 => n1901, B2 => n509, C1 => n1655, C2 => n510
                           , A => n511, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_24_port);
   U1957 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, A => n1706, ZN 
                           => n509);
   U1958 : AOI22_X1 port map( A1 => n1652, A2 => n512, B1 => 
                           DATAPATH_IxThird_stxALU1xN215, B2 => n1710, ZN => 
                           n511);
   U1959 : XNOR2_X1 port map( A => n471, B => n513, ZN => n510);
   U1960 : NAND2_X1 port map( A1 => n658, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, ZN => n647);
   U1961 : NAND2_X1 port map( A1 => n650, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n648);
   U1962 : NAND2_X1 port map( A1 => n605, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, ZN => n600);
   U1963 : NAND2_X1 port map( A1 => n695, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, ZN => n692);
   U1964 : OAI21_X1 port map( B1 => n783, B2 => n786, A => n600, ZN => n784);
   U1965 : NAND2_X1 port map( A1 => n601, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_16_port, ZN => n786);
   U1966 : AOI21_X1 port map( B1 => n1868, B2 => n1907, A => n555, ZN => n552);
   U1967 : INV_X1 port map( A => n543, ZN => n1907);
   U1968 : AOI21_X1 port map( B1 => n543, B2 => n520, A => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n555);
   U1969 : AOI21_X1 port map( B1 => n1864, B2 => n1902, A => n507, ZN => n504);
   U1970 : INV_X1 port map( A => n495, ZN => n1902);
   U1971 : AOI21_X1 port map( B1 => n495, B2 => n471, A => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, ZN => n507);
   U1972 : OAI221_X1 port map( B1 => n1910, B2 => n607, C1 => n1655, C2 => n608
                           , A => n609, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_17_port);
   U1973 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, A => n1706, ZN 
                           => n607);
   U1974 : AOI22_X1 port map( A1 => n1652, A2 => n610, B1 => 
                           DATAPATH_IxThird_stxALU1xN208, B2 => n1710, ZN => 
                           n609);
   U1975 : XNOR2_X1 port map( A => n611, B => n1871, ZN => n608);
   U1976 : OAI21_X1 port map( B1 => n171, B2 => n1646, A => n1767, ZN => n169);
   U1977 : AND2_X1 port map( A1 => n887, A2 => n1827, ZN => n870);
   U1978 : INV_X1 port map( A => n877, ZN => n1829);
   U1979 : INV_X1 port map( A => n165, ZN => n1851);
   U1980 : OAI21_X1 port map( B1 => n1608, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_12_port);
   U1981 : OAI21_X1 port map( B1 => n1609, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_13_port);
   U1982 : OAI21_X1 port map( B1 => n1615, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_14_port);
   U1983 : OAI21_X1 port map( B1 => n1624, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_29_port);
   U1984 : OAI21_X1 port map( B1 => n1386, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_31_port);
   U1985 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_18_port, ZN => 
                           n1870);
   U1986 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_10_port, ZN => 
                           n1879);
   U1987 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_14_port, ZN => 
                           n1875);
   U1988 : OAI21_X1 port map( B1 => n800, B2 => n801, A => n1964, ZN => n798);
   U1989 : BUF_X1 port map( A => n1635, Z => n1728);
   U1990 : INV_X1 port map( A => n878, ZN => n1825);
   U1991 : NOR2_X1 port map( A1 => n1646, A2 => n101, ZN => n106);
   U1992 : NAND2_X1 port map( A1 => n1826, A2 => n894, ZN => n874);
   U1993 : INV_X1 port map( A => n894, ZN => n1828);
   U1994 : INV_X1 port map( A => n872, ZN => n1827);
   U1995 : XNOR2_X1 port map( A => n814, B => n815, ZN => 
                           DATAPATH_IxSecond_stxjump_target_3_port);
   U1996 : NAND2_X1 port map( A1 => n1841, A2 => n284, ZN => n814);
   U1997 : INV_X1 port map( A => n817, ZN => n1841);
   U1998 : INV_X1 port map( A => n237, ZN => n1836);
   U1999 : INV_X1 port map( A => n1747, ZN => n1743);
   U2000 : XNOR2_X1 port map( A => n1663, B => n742, ZN => n495);
   U2001 : XNOR2_X1 port map( A => n1663, B => n750, ZN => n543);
   U2002 : INV_X1 port map( A => n109, ZN => n1767);
   U2003 : INV_X1 port map( A => n1732, ZN => n1731);
   U2004 : XNOR2_X1 port map( A => n1662, B => n735, ZN => n457);
   U2005 : OAI21_X1 port map( B1 => n1135, B2 => n1795, A => n1134, ZN => 
                           CU_IxN25);
   U2006 : INV_X1 port map( A => n27, ZN => n1795);
   U2007 : AOI21_X1 port map( B1 => n1137, B2 => n1797, A => n1138, ZN => n1135
                           );
   U2008 : XNOR2_X1 port map( A => n1661, B => n734, ZN => n729);
   U2009 : OAI221_X1 port map( B1 => n1654, B2 => n665, C1 => n1917, C2 => n667
                           , A => n668, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_11_port);
   U2010 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, A => n1705, ZN 
                           => n667);
   U2011 : AOI22_X1 port map( A1 => n1653, A2 => n669, B1 => 
                           DATAPATH_IxThird_stxALU1xN202, B2 => n1709, ZN => 
                           n668);
   U2012 : AOI22_X1 port map( A1 => n1882, A2 => n671, B1 => n672, B2 => n338, 
                           ZN => n665);
   U2013 : OAI221_X1 port map( B1 => n1655, B2 => n682, C1 => n1918, C2 => n684
                           , A => n685, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_10_port);
   U2014 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, A => n1705, ZN 
                           => n684);
   U2015 : AOI22_X1 port map( A1 => n1653, A2 => n686, B1 => 
                           DATAPATH_IxThird_stxALU1xN201, B2 => n1709, ZN => 
                           n685);
   U2016 : AOI22_X1 port map( A1 => n1882, A2 => n687, B1 => n688, B2 => n338, 
                           ZN => n682);
   U2017 : OAI221_X1 port map( B1 => n1654, B2 => n367, C1 => n1922, C2 => n369
                           , A => n370, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_6_port);
   U2018 : INV_X1 port map( A => n372, ZN => n1922);
   U2019 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_6_port, A => n1705, ZN 
                           => n369);
   U2020 : AOI22_X1 port map( A1 => n1651, A2 => n371, B1 => 
                           DATAPATH_IxThird_stxALU1xN197, B2 => n1711, ZN => 
                           n370);
   U2021 : OAI221_X1 port map( B1 => n1916, B2 => n660, C1 => n1655, C2 => n661
                           , A => n662, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_12_port);
   U2022 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, A => n1705, ZN 
                           => n660);
   U2023 : AOI22_X1 port map( A1 => n1653, A2 => n663, B1 => 
                           DATAPATH_IxThird_stxALU1xN203, B2 => n1709, ZN => 
                           n662);
   U2024 : XNOR2_X1 port map( A => n1877, B => n664, ZN => n661);
   U2025 : OAI221_X1 port map( B1 => n1919, B2 => n328, C1 => n1655, C2 => n330
                           , A => n331, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_9_port);
   U2026 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, A => n1705, ZN 
                           => n328);
   U2027 : AOI22_X1 port map( A1 => n1651, A2 => n333, B1 => 
                           DATAPATH_IxThird_stxALU1xN200, B2 => n1709, ZN => 
                           n331);
   U2028 : XNOR2_X1 port map( A => n335, B => n336, ZN => n330);
   U2029 : OAI221_X1 port map( B1 => n1732, B2 => n382, C1 => n1656, C2 => n383
                           , A => n384, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_5_port);
   U2030 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, A => n1705, ZN 
                           => n382);
   U2031 : AOI22_X1 port map( A1 => n1651, A2 => n385, B1 => 
                           DATAPATH_IxThird_stxALU1xN196, B2 => n1711, ZN => 
                           n384);
   U2032 : OAI221_X1 port map( B1 => n1734, B2 => n390, C1 => n1656, C2 => n391
                           , A => n392, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_4_port);
   U2033 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, A => n1705, ZN 
                           => n390);
   U2034 : AOI22_X1 port map( A1 => n1651, A2 => n393, B1 => 
                           DATAPATH_IxThird_stxALU1xN195, B2 => n1711, ZN => 
                           n392);
   U2035 : XNOR2_X1 port map( A => n394, B => n357, ZN => n391);
   U2036 : NOR2_X1 port map( A1 => n933, A2 => n941, ZN => n931);
   U2037 : XNOR2_X1 port map( A => n1668, B => n488, ZN => n481);
   U2038 : XNOR2_X1 port map( A => n1662, B => n741, ZN => n498);
   U2039 : XNOR2_X1 port map( A => n1664, B => n749, ZN => n546);
   U2040 : XNOR2_X1 port map( A => n1669, B => n747, ZN => n530);
   U2041 : NOR2_X1 port map( A1 => n605, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, ZN => n599);
   U2042 : NOR2_X1 port map( A1 => n498, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, ZN => n496);
   U2043 : NOR2_X1 port map( A1 => n546, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, ZN => n544);
   U2044 : NOR2_X1 port map( A1 => n695, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, ZN => n691);
   U2045 : NOR2_X1 port map( A1 => n457, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, ZN => n732);
   U2046 : NOR2_X1 port map( A1 => n650, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n646);
   U2047 : NOR2_X1 port map( A1 => n380, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, ZN => n377);
   U2048 : NOR2_X1 port map( A1 => n447, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, ZN => n443);
   U2049 : OAI221_X1 port map( B1 => n1654, B2 => n349, C1 => n1921, C2 => n351
                           , A => n352, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_7_port);
   U2050 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, A => n1705, ZN 
                           => n351);
   U2051 : AOI22_X1 port map( A1 => n1651, A2 => n353, B1 => 
                           DATAPATH_IxThird_stxALU1xN198, B2 => n1711, ZN => 
                           n352);
   U2052 : AOI22_X1 port map( A1 => n1886, A2 => n355, B1 => n356, B2 => n357, 
                           ZN => n349);
   U2053 : NOR2_X1 port map( A1 => n658, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, ZN => n649);
   U2054 : NOR2_X1 port map( A1 => n388, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, ZN => n376);
   U2055 : OAI21_X1 port map( B1 => n732, B2 => n1896, A => n733, ZN => n434);
   U2056 : OAI21_X1 port map( B1 => n729, B2 => n1857, A => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, ZN => n733);
   U2057 : OAI22_X1 port map( A1 => n1608, A2 => n1714, B1 => n1787, B2 => 
                           n1712, ZN => n1567);
   U2058 : OAI22_X1 port map( A1 => n1609, A2 => n1714, B1 => n1786, B2 => 
                           n1712, ZN => n1566);
   U2059 : OAI22_X1 port map( A1 => n1615, A2 => n1714, B1 => n1785, B2 => 
                           n1712, ZN => n1565);
   U2060 : OAI221_X1 port map( B1 => n1654, B2 => n620, C1 => n1913, C2 => n622
                           , A => n623, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_15_port);
   U2061 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_15_port, A => n1706, ZN 
                           => n622);
   U2062 : AOI22_X1 port map( A1 => n1653, A2 => n624, B1 => 
                           DATAPATH_IxThird_stxALU1xN206, B2 => n1709, ZN => 
                           n623);
   U2063 : AOI22_X1 port map( A1 => n625, A2 => n626, B1 => n1877, B2 => n628, 
                           ZN => n620);
   U2064 : OAI221_X1 port map( B1 => n1654, B2 => n638, C1 => n1914, C2 => n640
                           , A => n641, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_14_port);
   U2065 : AOI21_X1 port map( B1 => n1707, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_14_port, A => n1705, ZN 
                           => n640);
   U2066 : AOI22_X1 port map( A1 => n1653, A2 => n642, B1 => 
                           DATAPATH_IxThird_stxALU1xN205, B2 => n1709, ZN => 
                           n641);
   U2067 : AOI22_X1 port map( A1 => n643, A2 => n626, B1 => n1877, B2 => n644, 
                           ZN => n638);
   U2068 : OAI21_X1 port map( B1 => n1855, B2 => n1896, A => n728, ZN => n432);
   U2069 : OAI211_X1 port map( C1 => DATAPATH_IxThird_stxALU_IN1_29_port, C2 =>
                           n729, A => DATAPATH_IxThird_stxALU_IN1_28_port, B =>
                           n457, ZN => n728);
   U2070 : OAI21_X1 port map( B1 => n497, B2 => n496, A => n492, ZN => n480);
   U2071 : NOR2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_24_port, A2 => 
                           n495, ZN => n497);
   U2072 : OAI21_X1 port map( B1 => n545, B2 => n544, A => n540, ZN => n529);
   U2073 : NOR2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_20_port, A2 => 
                           n543, ZN => n545);
   U2074 : OAI21_X1 port map( B1 => n598, B2 => n599, A => n600, ZN => n583);
   U2075 : NOR2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_16_port, A2 => 
                           n601, ZN => n598);
   U2076 : INV_X1 port map( A => CU_IxN24, ZN => n1753);
   U2077 : OAI221_X1 port map( B1 => n1920, B2 => n344, C1 => n1656, C2 => n345
                           , A => n346, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_8_port);
   U2078 : AOI21_X1 port map( B1 => n1708, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, A => n1705, ZN 
                           => n344);
   U2079 : AOI22_X1 port map( A1 => n1651, A2 => n347, B1 => 
                           DATAPATH_IxThird_stxALU1xN199, B2 => n1711, ZN => 
                           n346);
   U2080 : XNOR2_X1 port map( A => n338, B => n348, ZN => n345);
   U2081 : NOR2_X1 port map( A1 => n569, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_0_port, ZN => n442);
   U2082 : NAND2_X1 port map( A1 => n498, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, ZN => n492);
   U2083 : NAND2_X1 port map( A1 => n546, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, ZN => n540);
   U2084 : XNOR2_X1 port map( A => n1337, B => n731, ZN => n730);
   U2085 : OAI21_X1 port map( B1 => n690, B2 => n691, A => n692, ZN => n675);
   U2086 : NOR2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_8_port, A2 => 
                           n337, ZN => n690);
   U2087 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_2_port, Z => n1738
                           );
   U2088 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_3_port, Z => n1736
                           );
   U2089 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_16_port, ZN => 
                           n1872);
   U2090 : NOR2_X1 port map( A1 => CU_Ixcw_LUT_16_port, A2 => n326, ZN => 
                           CU_Ixcw1_14_port);
   U2091 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_29_port, ZN => 
                           n1855);
   U2092 : INV_X1 port map( A => n91, ZN => n1757);
   U2093 : OAI21_X1 port map( B1 => CU_Ixcw_LUT_15_port, B2 => n1746, A => 
                           n1716, ZN => n91);
   U2094 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_0_port, Z => n1742
                           );
   U2095 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_1_port, Z => n1740
                           );
   U2096 : NAND2_X1 port map( A1 => n326, A2 => n1743, ZN => n92);
   U2097 : INV_X1 port map( A => n159, ZN => n1852);
   U2098 : BUF_X1 port map( A => n1635, Z => n1727);
   U2099 : BUF_X1 port map( A => n1635, Z => n1726);
   U2100 : BUF_X1 port map( A => n1635, Z => n1725);
   U2101 : BUF_X1 port map( A => n1635, Z => n1724);
   U2102 : BUF_X1 port map( A => n1635, Z => n1723);
   U2103 : BUF_X1 port map( A => n1635, Z => n1722);
   U2104 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_22_port, ZN => 
                           n1866);
   U2105 : AND2_X1 port map( A1 => n730, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, ZN => n719);
   U2106 : BUF_X1 port map( A => n1621, Z => n1658);
   U2107 : INV_X1 port map( A => n171, ZN => n1971);
   U2108 : INV_X1 port map( A => n1138, ZN => n1794);
   U2109 : INV_X1 port map( A => n256, ZN => n1977);
   U2110 : INV_X1 port map( A => n224, ZN => n1974);
   U2111 : INV_X1 port map( A => n234, ZN => n1975);
   U2112 : INV_X1 port map( A => n246, ZN => n1976);
   U2113 : INV_X1 port map( A => n214, ZN => n1973);
   U2114 : INV_X1 port map( A => n192, ZN => n1972);
   U2115 : NAND2_X1 port map( A1 => n492, A2 => n493, ZN => n476);
   U2116 : INV_X1 port map( A => n496, ZN => n1863);
   U2117 : NAND2_X1 port map( A1 => n540, A2 => n541, ZN => n525);
   U2118 : INV_X1 port map( A => n544, ZN => n1867);
   U2119 : NAND2_X1 port map( A1 => n692, A2 => n693, ZN => n679);
   U2120 : INV_X1 port map( A => n691, ZN => n1880);
   U2121 : INV_X1 port map( A => n789, ZN => n1898);
   U2122 : INV_X1 port map( A => n118, ZN => n1970);
   U2123 : NAND2_X1 port map( A1 => n1965, A2 => n809, ZN => n813);
   U2124 : OR2_X1 port map( A1 => n730, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, ZN => n727);
   U2125 : AND2_X1 port map( A1 => n1767, A2 => n289, ZN => n285);
   U2126 : INV_X1 port map( A => n298, ZN => n1924);
   U2127 : INV_X1 port map( A => n811, ZN => n1965);
   U2128 : INV_X1 port map( A => CU_IxN23, ZN => n1752);
   U2129 : OAI21_X1 port map( B1 => n337, B2 => n338, A => n1881, ZN => n335);
   U2130 : INV_X1 port map( A => n340, ZN => n1881);
   U2131 : AOI21_X1 port map( B1 => n338, B2 => n337, A => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, ZN => n340);
   U2132 : INV_X1 port map( A => n949, ZN => n1962);
   U2133 : AND2_X1 port map( A1 => CU_Ixcw_LUT_0_port, A2 => n1853, ZN => 
                           CU_Ixcw1_0_port);
   U2134 : AND2_X1 port map( A1 => CU_Ixcw_LUT_8_port, A2 => n1853, ZN => 
                           CU_Ixcw1_8_port);
   U2135 : AND2_X1 port map( A1 => CU_Ixcw_LUT_4_port, A2 => n1853, ZN => 
                           CU_Ixcw1_4_port);
   U2136 : AND2_X1 port map( A1 => CU_Ixcw_LUT_2_port, A2 => n1853, ZN => 
                           CU_Ixcw1_2_port);
   U2137 : AND2_X1 port map( A1 => CU_Ixcw_LUT_1_port, A2 => n1853, ZN => 
                           CU_Ixcw1_1_port);
   U2138 : AND2_X1 port map( A1 => CU_Ixcw_LUT_5_port, A2 => n1853, ZN => 
                           CU_Ixcw1_5_port);
   U2139 : AND2_X1 port map( A1 => CU_Ixcw_LUT_7_port, A2 => n1853, ZN => 
                           CU_Ixcw1_7_port);
   U2140 : NOR3_X1 port map( A1 => n1794, A2 => n1745, A3 => n1797, ZN => n28);
   U2141 : AOI21_X1 port map( B1 => n1618, B2 => n1659, A => n843, ZN => n834);
   U2142 : AOI21_X1 port map( B1 => n1619, B2 => n1658, A => n860, ZN => n851);
   U2143 : BUF_X1 port map( A => n334, Z => n1709);
   U2144 : INV_X1 port map( A => n1636, ZN => n1707);
   U2145 : BUF_X1 port map( A => n334, Z => n1710);
   U2146 : INV_X1 port map( A => n1636, ZN => n1708);
   U2147 : OAI21_X1 port map( B1 => n1672, B2 => n1591, A => n790, ZN => n421);
   U2148 : BUF_X1 port map( A => n334, Z => n1711);
   U2149 : OAI21_X1 port map( B1 => n949, B2 => n794, A => n950, ZN => n942);
   U2150 : INV_X1 port map( A => n570, ZN => n1890);
   U2151 : AOI21_X1 port map( B1 => DATAPATH_IxThird_stxALU_IN1_1_port, B2 => 
                           n1707, A => n1706, ZN => n570);
   U2152 : INV_X1 port map( A => n705, ZN => n1891);
   U2153 : AOI21_X1 port map( B1 => DATAPATH_IxThird_stxALU_IN1_0_port, B2 => 
                           n1707, A => n1706, ZN => n705);
   U2154 : AOI21_X1 port map( B1 => n1659, B2 => n1617, A => n824, ZN => n821);
   U2155 : OAI21_X1 port map( B1 => n1887, B2 => n1636, A => n1590, ZN => n400)
                           ;
   U2156 : OAI21_X1 port map( B1 => n1889, B2 => n1636, A => n1590, ZN => n439)
                           ;
   U2157 : BUF_X1 port map( A => n1621, Z => n1659);
   U2158 : OAI21_X1 port map( B1 => n1660, B2 => n1617, A => n826, ZN => n825);
   U2159 : INV_X1 port map( A => n418, ZN => n1925);
   U2160 : OAI21_X1 port map( B1 => n941, B2 => n946, A => n1961, ZN => n944);
   U2161 : BUF_X1 port map( A => n1657, Z => n1660);
   U2162 : BUF_X1 port map( A => n1659, Z => n1657);
   U2163 : INV_X1 port map( A => n933, ZN => n1961);
   U2164 : INV_X1 port map( A => n805, ZN => n1964);
   U2165 : AOI22_X1 port map( A1 => RF_WR_DATAx24x, A2 => n1698, B1 => 
                           RF_RD1_DATA(24), B2 => n1695, ZN => n1019);
   U2166 : AOI22_X1 port map( A1 => RF_WR_DATAx20x, A2 => n1697, B1 => 
                           RF_RD1_DATA(20), B2 => n1696, ZN => n994);
   U2167 : AOI22_X1 port map( A1 => RF_WR_DATAx8x, A2 => n1698, B1 => 
                           RF_RD1_DATA(8), B2 => n1695, ZN => n1037);
   U2168 : AOI22_X1 port map( A1 => RF_WR_DATAx28x, A2 => n1698, B1 => 
                           RF_RD1_DATA(28), B2 => n1695, ZN => n1029);
   U2169 : AOI22_X1 port map( A1 => RF_WR_DATAx16x, A2 => n1697, B1 => 
                           RF_RD1_DATA(16), B2 => n1696, ZN => n991);
   U2170 : AOI22_X1 port map( A1 => RF_RD1_DATA(29), A2 => n1694, B1 => 
                           RF_WR_DATAx29x, B2 => n1697, ZN => n1032);
   U2171 : OAI221_X1 port map( B1 => n1702, B2 => n1583, C1 => n1440, C2 => 
                           n1699, A => n997, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_21_port);
   U2172 : AOI22_X1 port map( A1 => RF_WR_DATAx21x, A2 => n1697, B1 => 
                           RF_RD1_DATA(21), B2 => n1696, ZN => n997);
   U2173 : OAI221_X1 port map( B1 => n1703, B2 => n1594, C1 => n1428, C2 => 
                           n1700, A => n1040, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_9_port);
   U2174 : AOI22_X1 port map( A1 => RF_WR_DATAx9x, A2 => n1698, B1 => 
                           RF_RD1_DATA(9), B2 => n1695, ZN => n1040);
   U2175 : OAI221_X1 port map( B1 => n1702, B2 => n1604, C1 => n1436, C2 => 
                           n1699, A => n1007, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_17_port);
   U2176 : AOI22_X1 port map( A1 => RF_WR_DATAx17x, A2 => n1697, B1 => 
                           RF_RD1_DATA(17), B2 => n1696, ZN => n1007);
   U2177 : OAI22_X1 port map( A1 => n1353, A2 => n867, B1 => n868, B2 => n869, 
                           ZN => n181);
   U2178 : AOI21_X1 port map( B1 => n870, B2 => n871, A => n872, ZN => n868);
   U2179 : OAI21_X1 port map( B1 => n873, B2 => n874, A => n1826, ZN => n871);
   U2180 : AOI21_X1 port map( B1 => n876, B2 => n877, A => n878, ZN => n873);
   U2181 : NOR2_X2 port map( A1 => n1853, A2 => n1298, ZN => n291);
   U2182 : OAI221_X1 port map( B1 => n1704, B2 => n1599, C1 => n1420, C2 => 
                           n1701, A => n1086, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_1_port);
   U2183 : AOI22_X1 port map( A1 => RF_WR_DATAx1x, A2 => n1698, B1 => 
                           RF_RD1_DATA(1), B2 => n1695, ZN => n1086);
   U2184 : OAI221_X1 port map( B1 => n1702, B2 => n1584, C1 => n1449, C2 => 
                           n1699, A => n1010, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_30_port);
   U2185 : AOI22_X1 port map( A1 => RF_WR_DATAx30x, A2 => n1698, B1 => 
                           RF_RD1_DATA(30), B2 => n1696, ZN => n1010);
   U2186 : OAI221_X1 port map( B1 => n1702, B2 => n1588, C1 => n1442, C2 => 
                           n1699, A => n1000, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_23_port);
   U2187 : AOI22_X1 port map( A1 => RF_WR_DATAx23x, A2 => n1697, B1 => 
                           RF_RD1_DATA(23), B2 => n1696, ZN => n1000);
   U2188 : OAI221_X1 port map( B1 => n1702, B2 => n1586, C1 => n1441, C2 => 
                           n1699, A => n988, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_22_port);
   U2189 : AOI22_X1 port map( A1 => RF_WR_DATAx22x, A2 => n1697, B1 => 
                           RF_RD1_DATA(22), B2 => n1696, ZN => n988);
   U2190 : OAI221_X1 port map( B1 => n1702, B2 => n1600, C1 => n1438, C2 => 
                           n1699, A => n977, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_19_port);
   U2191 : AOI22_X1 port map( A1 => RF_WR_DATAx19x, A2 => n1697, B1 => 
                           RF_RD1_DATA(19), B2 => n1694, ZN => n977);
   U2192 : OAI221_X1 port map( B1 => n1703, B2 => n1601, C1 => n1430, C2 => 
                           n1700, A => n1057, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_11_port);
   U2193 : AOI22_X1 port map( A1 => RF_WR_DATAx11x, A2 => n1697, B1 => 
                           RF_RD1_DATA(11), B2 => n1695, ZN => n1057);
   U2194 : OAI221_X1 port map( B1 => n1704, B2 => n1578, C1 => n1426, C2 => 
                           n1701, A => n1064, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_7_port);
   U2195 : AOI22_X1 port map( A1 => RF_WR_DATAx7x, A2 => n1697, B1 => 
                           RF_RD1_DATA(7), B2 => n1694, ZN => n1064);
   U2196 : OAI221_X1 port map( B1 => n1702, B2 => n1603, C1 => n1437, C2 => 
                           n1699, A => n1004, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_18_port);
   U2197 : AOI22_X1 port map( A1 => RF_WR_DATAx18x, A2 => n1698, B1 => 
                           RF_RD1_DATA(18), B2 => n1696, ZN => n1004);
   U2198 : OAI221_X1 port map( B1 => n1703, B2 => n1607, C1 => n1429, C2 => 
                           n1700, A => n1054, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_10_port);
   U2199 : AOI22_X1 port map( A1 => RF_WR_DATAx10x, A2 => n1697, B1 => 
                           RF_RD1_DATA(10), B2 => n1694, ZN => n1054);
   U2200 : AOI211_X1 port map( C1 => n1608, C2 => n1830, A => n896, B => n1347,
                           ZN => n921);
   U2201 : AOI211_X1 port map( C1 => n1615, C2 => n1830, A => n896, B => n1349,
                           ZN => n907);
   U2202 : AOI211_X1 port map( C1 => n1609, C2 => n1830, A => n896, B => n1348,
                           ZN => n922);
   U2203 : OAI22_X1 port map( A1 => n1346, A2 => n1833, B1 => n929, B2 => n930,
                           ZN => n919);
   U2204 : AOI21_X1 port map( B1 => n931, B2 => n932, A => n933, ZN => n929);
   U2205 : OAI21_X1 port map( B1 => n934, B2 => n791, A => n1962, ZN => n932);
   U2206 : AOI21_X1 port map( B1 => n244, B2 => n936, A => n794, ZN => n934);
   U2207 : OAI221_X1 port map( B1 => n1425, B2 => n1693, C1 => n1190, C2 => 
                           n1690, A => n1078, ZN => n372);
   U2208 : AOI22_X1 port map( A1 => RF_WR_DATAx6x, A2 => n1686, B1 => 
                           RF_RD2_DATA(6), B2 => n1685, ZN => n1078);
   U2209 : OAI221_X1 port map( B1 => n1445, B2 => n1692, C1 => n1168, C2 => 
                           n1689, A => n1024, ZN => n488);
   U2210 : AOI22_X1 port map( A1 => RF_WR_DATAx26x, A2 => n1687, B1 => 
                           RF_RD2_DATA(26), B2 => n1684, ZN => n1024);
   U2211 : OAI22_X1 port map( A1 => n1383, A2 => n1611, B1 => n952, B2 => n799,
                           ZN => n936);
   U2212 : AOI21_X1 port map( B1 => n808, B2 => n953, A => n805, ZN => n952);
   U2213 : OAI21_X1 port map( B1 => n954, B2 => n813, A => n1965, ZN => n953);
   U2214 : AOI21_X1 port map( B1 => n1844, B2 => n1838, A => n270, ZN => n954);
   U2215 : OAI211_X1 port map( C1 => n1357, C2 => n1386, A => n850, B => n851, 
                           ZN => n835);
   U2216 : NAND4_X1 port map( A1 => n180, A2 => n181, A3 => n852, A4 => n853, 
                           ZN => n850);
   U2217 : NOR2_X1 port map( A1 => n854, A2 => n855, ZN => n853);
   U2218 : OAI221_X1 port map( B1 => n1704, B2 => n1595, C1 => n1425, C2 => 
                           n1701, A => n1077, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_6_port);
   U2219 : AOI22_X1 port map( A1 => RF_WR_DATAx6x, A2 => n1697, B1 => 
                           RF_RD1_DATA(6), B2 => n1694, ZN => n1077);
   U2220 : OAI221_X1 port map( B1 => n1703, B2 => n1585, C1 => n1445, C2 => 
                           n1700, A => n1023, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_26_port);
   U2221 : AOI22_X1 port map( A1 => RF_WR_DATAx26x, A2 => n1698, B1 => 
                           RF_RD1_DATA(26), B2 => n1695, ZN => n1023);
   U2222 : NAND2_X1 port map( A1 => CU_Ixcw2_i_12_port, A2 => n1850, ZN => n897
                           );
   U2223 : OAI221_X1 port map( B1 => n1440, B2 => n1691, C1 => n1173, C2 => 
                           n1688, A => n998, ZN => n749);
   U2224 : AOI22_X1 port map( A1 => RF_WR_DATAx21x, A2 => n1687, B1 => 
                           RF_RD2_DATA(21), B2 => n1683, ZN => n998);
   U2225 : OAI221_X1 port map( B1 => n1449, B2 => n1691, C1 => n1169, C2 => 
                           n1688, A => n1011, ZN => n731);
   U2226 : AOI22_X1 port map( A1 => RF_WR_DATAx30x, A2 => n1687, B1 => 
                           RF_RD2_DATA(30), B2 => n1683, ZN => n1011);
   U2227 : OAI221_X1 port map( B1 => n1436, B2 => n1691, C1 => n1176, C2 => 
                           n1688, A => n1008, ZN => n787);
   U2228 : AOI22_X1 port map( A1 => RF_WR_DATAx17x, A2 => n1687, B1 => 
                           RF_RD2_DATA(17), B2 => n1683, ZN => n1008);
   U2229 : OAI221_X1 port map( B1 => n1448, B2 => n1692, C1 => n1157, C2 => 
                           n1689, A => n1033, ZN => n734);
   U2230 : AOI22_X1 port map( A1 => RF_WR_DATAx29x, A2 => n1687, B1 => 
                           RF_RD2_DATA(29), B2 => n1684, ZN => n1033);
   U2231 : OAI221_X1 port map( B1 => n1435, B2 => n1691, C1 => n1180, C2 => 
                           n1688, A => n992, ZN => n788);
   U2232 : AOI22_X1 port map( A1 => RF_WR_DATAx16x, A2 => n1686, B1 => 
                           RF_RD2_DATA(16), B2 => n1683, ZN => n992);
   U2233 : OAI221_X1 port map( B1 => n1427, B2 => n1692, C1 => n1185, C2 => 
                           n1689, A => n1038, ZN => n771);
   U2234 : AOI22_X1 port map( A1 => RF_WR_DATAx8x, A2 => n1687, B1 => 
                           RF_RD2_DATA(8), B2 => n1684, ZN => n1038);
   U2235 : OAI221_X1 port map( B1 => n1439, B2 => n1691, C1 => n1178, C2 => 
                           n1688, A => n995, ZN => n750);
   U2236 : AOI22_X1 port map( A1 => RF_WR_DATAx20x, A2 => n1686, B1 => 
                           RF_RD2_DATA(20), B2 => n1683, ZN => n995);
   U2237 : OAI221_X1 port map( B1 => n1432, B2 => n1692, C1 => n1188, C2 => 
                           n1689, A => n1062, ZN => n762);
   U2238 : AOI22_X1 port map( A1 => RF_WR_DATAx13x, A2 => n1686, B1 => 
                           RF_RD2_DATA(13), B2 => n1684, ZN => n1062);
   U2239 : OAI221_X1 port map( B1 => n1437, B2 => n1691, C1 => n1175, C2 => 
                           n1688, A => n1005, ZN => n785);
   U2240 : AOI22_X1 port map( A1 => RF_WR_DATAx18x, A2 => n1687, B1 => 
                           RF_RD2_DATA(18), B2 => n1683, ZN => n1005);
   U2241 : OAI221_X1 port map( B1 => n1441, B2 => n1691, C1 => n1179, C2 => 
                           n1688, A => n989, ZN => n747);
   U2242 : AOI22_X1 port map( A1 => RF_WR_DATAx22x, A2 => n1686, B1 => 
                           RF_RD2_DATA(22), B2 => n1683, ZN => n989);
   U2243 : OAI221_X1 port map( B1 => n1433, B2 => n1692, C1 => n1183, C2 => 
                           n1689, A => n1044, ZN => n760);
   U2244 : AOI22_X1 port map( A1 => RF_WR_DATAx14x, A2 => n1687, B1 => 
                           RF_RD2_DATA(14), B2 => n1684, ZN => n1044);
   U2245 : OAI221_X1 port map( B1 => n1446, B2 => n1692, C1 => n1167, C2 => 
                           n1689, A => n1027, ZN => n789);
   U2246 : AOI22_X1 port map( A1 => RF_WR_DATAx27x, A2 => n1687, B1 => 
                           RF_RD2_DATA(27), B2 => n1684, ZN => n1027);
   U2247 : OAI211_X1 port map( C1 => n897, C2 => n1608, A => n1830, B => n1347,
                           ZN => n912);
   U2248 : OAI211_X1 port map( C1 => n1361, C2 => n1386, A => n833, B => n834, 
                           ZN => n819);
   U2249 : NAND4_X1 port map( A1 => n152, A2 => n835, A3 => n836, A4 => n837, 
                           ZN => n833);
   U2250 : NOR2_X1 port map( A1 => n838, A2 => n839, ZN => n837);
   U2251 : OAI211_X1 port map( C1 => n897, C2 => n1609, A => n1830, B => n1348,
                           ZN => n911);
   U2252 : XNOR2_X1 port map( A => n1362, B => n1657, ZN => n126);
   U2253 : OAI221_X1 port map( B1 => n1419, B2 => n1693, C1 => n1193, C2 => 
                           n1690, A => n1069, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_0_port);
   U2254 : AOI22_X1 port map( A1 => RF_WR_DATAx0x, A2 => n1686, B1 => 
                           RF_RD2_DATA(0), B2 => n1685, ZN => n1069);
   U2255 : OAI221_X1 port map( B1 => n1420, B2 => n1693, C1 => n1194, C2 => 
                           n1690, A => n1109, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_1_port);
   U2256 : AOI22_X1 port map( A1 => RF_WR_DATAx1x, A2 => n1687, B1 => 
                           RF_RD2_DATA(1), B2 => n1685, ZN => n1109);
   U2257 : OAI221_X1 port map( B1 => n1421, B2 => n1693, C1 => n1195, C2 => 
                           n1690, A => n1081, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_2_port);
   U2258 : AOI22_X1 port map( A1 => n1687, A2 => RF_WR_DATAx2x, B1 => 
                           RF_RD2_DATA(2), B2 => n1685, ZN => n1081);
   U2259 : OAI221_X1 port map( B1 => n1422, B2 => n1693, C1 => n1196, C2 => 
                           n1690, A => n1084, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_3_port);
   U2260 : AOI22_X1 port map( A1 => RF_WR_DATAx3x, A2 => n1686, B1 => 
                           RF_RD2_DATA(3), B2 => n1685, ZN => n1084);
   U2261 : NOR4_X1 port map( A1 => n971, A2 => n972, A3 => n973, A4 => n974, ZN
                           => n970);
   U2262 : NAND4_X1 port map( A1 => n1856, A2 => BRANCH_EN_i, A3 => n463, A4 =>
                           n1022, ZN => n971);
   U2263 : OR4_X1 port map( A1 => n610, A2 => n594, A3 => n518, A4 => n551, ZN 
                           => n973);
   U2264 : OR4_X1 port map( A1 => n560, A2 => n618, A3 => n536, A4 => n576, ZN 
                           => n974);
   U2265 : NOR4_X1 port map( A1 => n1299, A2 => n1120, A3 => n1130, A4 => n1131
                           , ZN => n1129);
   U2266 : NOR4_X1 port map( A1 => n1299, A2 => n1096, A3 => n1106, A4 => n1107
                           , ZN => n1105);
   U2267 : OAI221_X1 port map( B1 => n1450, B2 => n1691, C1 => n1170, C2 => 
                           n1688, A => n1014, ZN => n715);
   U2268 : AOI22_X1 port map( A1 => RF_WR_DATAx31x, A2 => n1687, B1 => 
                           RF_RD2_DATA(31), B2 => n1683, ZN => n1014);
   U2269 : AOI21_X1 port map( B1 => n1614, B2 => n958, A => n959, ZN => n268);
   U2270 : AOI21_X1 port map( B1 => n282, B2 => n284, A => n815, ZN => n959);
   U2271 : NAND2_X1 port map( A1 => n1118, A2 => n1119, ZN => n1116);
   U2272 : NOR4_X1 port map( A1 => n1122, A2 => n1123, A3 => n1124, A4 => n1125
                           , ZN => n1118);
   U2273 : NOR4_X1 port map( A1 => n1333, A2 => n1334, A3 => n1120, A4 => n1121
                           , ZN => n1119);
   U2274 : NAND2_X1 port map( A1 => n1094, A2 => n1095, ZN => n1092);
   U2275 : NOR4_X1 port map( A1 => n1098, A2 => n1099, A3 => n1100, A4 => n1101
                           , ZN => n1094);
   U2276 : NOR4_X1 port map( A1 => n1333, A2 => n1334, A3 => n1096, A4 => n1097
                           , ZN => n1095);
   U2277 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_5_port, ZN => 
                           n1732);
   U2278 : OAI221_X1 port map( B1 => n1424, B2 => n1693, C1 => n1191, C2 => 
                           n1690, A => n1075, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_5_port);
   U2279 : AOI22_X1 port map( A1 => RF_WR_DATAx5x, A2 => n1686, B1 => 
                           RF_RD2_DATA(5), B2 => n1685, ZN => n1075);
   U2280 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_4_port, ZN => 
                           n1734);
   U2281 : OAI221_X1 port map( B1 => n1423, B2 => n1693, C1 => n1192, C2 => 
                           n1690, A => n1072, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_4_port);
   U2282 : AOI22_X1 port map( A1 => RF_WR_DATAx4x, A2 => n1686, B1 => 
                           RF_RD2_DATA(4), B2 => n1685, ZN => n1072);
   U2283 : OAI221_X1 port map( B1 => n1704, B2 => n1579, C1 => n1421, C2 => 
                           n1701, A => n1080, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_2_port);
   U2284 : AOI22_X1 port map( A1 => n1697, A2 => RF_WR_DATAx2x, B1 => 
                           RF_RD1_DATA(2), B2 => n1694, ZN => n1080);
   U2285 : OAI221_X1 port map( B1 => n1704, B2 => n1597, C1 => n1422, C2 => 
                           n1701, A => n1083, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_3_port);
   U2286 : AOI22_X1 port map( A1 => RF_WR_DATAx3x, A2 => n1697, B1 => 
                           RF_RD1_DATA(3), B2 => n1694, ZN => n1083);
   U2287 : AOI22_X1 port map( A1 => n897, A2 => n1368, B1 => n1847, B2 => n1378
                           , ZN => n283);
   U2288 : AOI21_X1 port map( B1 => n294, B2 => n298, A => n1197, ZN => n326);
   U2289 : OAI22_X1 port map( A1 => n1409, A2 => n1767, B1 => n109, B2 => n158,
                           ZN => n1525);
   U2290 : AOI211_X1 port map( C1 => n159, C2 => 
                           DATAPATH_IxSecond_stxjump_target_22_port, A => n160,
                           B => n161, ZN => n158);
   U2291 : OAI21_X1 port map( B1 => n1228, B2 => n165, A => n1743, ZN => n160);
   U2292 : NOR3_X1 port map( A1 => n162, A2 => n1851, A3 => n159, ZN => n161);
   U2293 : INV_X1 port map( A => n1065, ZN => n1921);
   U2294 : OAI221_X1 port map( B1 => n1426, B2 => n1693, C1 => n1189, C2 => 
                           n1690, A => n1066, ZN => n1065);
   U2295 : AOI22_X1 port map( A1 => RF_WR_DATAx7x, A2 => n1686, B1 => 
                           RF_RD2_DATA(7), B2 => n1685, ZN => n1066);
   U2296 : OAI22_X1 port map( A1 => n1370, A2 => n1847, B1 => n1380, B2 => n897
                           , ZN => n956);
   U2297 : OAI22_X1 port map( A1 => n1815, A2 => n818, B1 => n819, B2 => n820, 
                           ZN => DATAPATH_IxSecond_stxjump_target_31_port);
   U2298 : OAI22_X1 port map( A1 => n1815, A2 => n827, B1 => n828, B2 => n819, 
                           ZN => DATAPATH_IxSecond_stxjump_target_30_port);
   U2299 : XNOR2_X1 port map( A => n1364, B => n1386, ZN => n829);
   U2300 : AOI22_X1 port map( A1 => n897, A2 => n1367, B1 => n1847, B2 => n1377
                           , ZN => n286);
   U2301 : XNOR2_X1 port map( A => n1833, B => n1346, ZN => n930);
   U2302 : AOI21_X1 port map( B1 => n1830, B2 => n1371, A => n896, ZN => n913);
   U2303 : AOI22_X1 port map( A1 => n897, A2 => n1369, B1 => n1847, B2 => n1379
                           , ZN => n958);
   U2304 : OAI21_X1 port map( B1 => n1967, B2 => IMM_SEL_i, A => n1116, ZN => 
                           n1111);
   U2305 : INV_X1 port map( A => n1115, ZN => n1967);
   U2306 : OAI21_X1 port map( B1 => n1969, B2 => PC_SEL_i, A => n1092, ZN => 
                           n1088);
   U2307 : INV_X1 port map( A => n1093, ZN => n1969);
   U2308 : OAI221_X1 port map( B1 => n1235, B2 => n1649, C1 => n111, C2 => 
                           n1647, A => n112, ZN => n1518);
   U2309 : AOI21_X1 port map( B1 => n113, B2 => IRAM_ADD_29_port, A => n115, ZN
                           => n112);
   U2310 : NOR3_X1 port map( A1 => IRAM_ADD_29_port, A2 => n110, A3 => n1644, 
                           ZN => n115);
   U2311 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_28_port, A => n119, 
                           ZN => n113);
   U2312 : OAI221_X1 port map( B1 => n1647, B2 => n47, C1 => n1234, C2 => n1649
                           , A => n120, ZN => n1519);
   U2313 : AOI21_X1 port map( B1 => n1758, B2 => IRAM_ADD_28_port, A => n122, 
                           ZN => n120);
   U2314 : NOR4_X1 port map( A1 => n1414, A2 => n1970, A3 => n1644, A4 => 
                           IRAM_ADD_28_port, ZN => n122);
   U2315 : INV_X1 port map( A => n119, ZN => n1758);
   U2316 : OAI221_X1 port map( B1 => n1233, B2 => n1649, C1 => n1807, C2 => 
                           n1647, A => n129, ZN => n1520);
   U2317 : AOI21_X1 port map( B1 => n124, B2 => IRAM_ADD_27_port, A => n130, ZN
                           => n129);
   U2318 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_27_port, ZN 
                           => n1807);
   U2319 : NOR3_X1 port map( A1 => IRAM_ADD_27_port, A2 => n1970, A3 => n1644, 
                           ZN => n130);
   U2320 : OAI221_X1 port map( B1 => n1232, B2 => n1649, C1 => n1808, C2 => 
                           n1647, A => n134, ZN => n1521);
   U2321 : AOI21_X1 port map( B1 => n135, B2 => IRAM_ADD_26_port, A => n137, ZN
                           => n134);
   U2322 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_26_port, ZN 
                           => n1808);
   U2323 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_25_port, A => n139, 
                           ZN => n135);
   U2324 : OAI221_X1 port map( B1 => n1231, B2 => n1649, C1 => n1809, C2 => 
                           n1647, A => n141, ZN => n1522);
   U2325 : AOI21_X1 port map( B1 => n1763, B2 => IRAM_ADD_25_port, A => n143, 
                           ZN => n141);
   U2326 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_25_port, ZN 
                           => n1809);
   U2327 : INV_X1 port map( A => n139, ZN => n1763);
   U2328 : OAI221_X1 port map( B1 => n1647, B2 => n46, C1 => n1230, C2 => n1649
                           , A => n145, ZN => n1523);
   U2329 : AOI21_X1 port map( B1 => n146, B2 => IRAM_ADD_24_port, A => n148, ZN
                           => n145);
   U2330 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_23_port, A => n150, 
                           ZN => n146);
   U2331 : NOR4_X1 port map( A1 => n1410, A2 => n144, A3 => n1644, A4 => 
                           IRAM_ADD_24_port, ZN => n148);
   U2332 : OAI221_X1 port map( B1 => n1229, B2 => n1649, C1 => n1803, C2 => 
                           n1647, A => n154, ZN => n1524);
   U2333 : AOI21_X1 port map( B1 => n1762, B2 => IRAM_ADD_23_port, A => n156, 
                           ZN => n154);
   U2334 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_23_port, ZN 
                           => n1803);
   U2335 : INV_X1 port map( A => n150, ZN => n1762);
   U2336 : OAI221_X1 port map( B1 => n1227, B2 => n1649, C1 => n1804, C2 => 
                           n1647, A => n167, ZN => n1526);
   U2337 : AOI22_X1 port map( A1 => n168, A2 => n1408, B1 => n169, B2 => 
                           IRAM_ADD_21_port, ZN => n167);
   U2338 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_21_port, ZN 
                           => n1804);
   U2339 : OAI221_X1 port map( B1 => n1225, B2 => n1649, C1 => n1648, C2 => 
                           n182, A => n183, ZN => n1528);
   U2340 : AOI21_X1 port map( B1 => n1761, B2 => IRAM_ADD_19_port, A => n185, 
                           ZN => n183);
   U2341 : INV_X1 port map( A => n179, ZN => n1761);
   U2342 : NOR3_X1 port map( A1 => IRAM_ADD_19_port, A2 => n172, A3 => n1645, 
                           ZN => n185);
   U2343 : OAI221_X1 port map( B1 => n1224, B2 => n1650, C1 => n1818, C2 => 
                           n1647, A => n196, ZN => n1530);
   U2344 : AOI21_X1 port map( B1 => n194, B2 => IRAM_ADD_17_port, A => n197, ZN
                           => n196);
   U2345 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_17_port, ZN 
                           => n1818);
   U2346 : NOR3_X1 port map( A1 => IRAM_ADD_17_port, A2 => n1972, A3 => n1645, 
                           ZN => n197);
   U2347 : OAI221_X1 port map( B1 => n1223, B2 => n1650, C1 => n1817, C2 => 
                           n1648, A => n200, ZN => n1531);
   U2348 : AOI21_X1 port map( B1 => n201, B2 => IRAM_ADD_16_port, A => n203, ZN
                           => n200);
   U2349 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_16_port, ZN 
                           => n1817);
   U2350 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_15_port, A => n205, 
                           ZN => n201);
   U2351 : XNOR2_X1 port map( A => n913, B => n1257, ZN => n904);
   U2352 : AOI211_X1 port map( C1 => n1860, C2 => n706, A => n1335, B => n1664,
                           ZN => n703);
   U2353 : OAI221_X1 port map( B1 => n1444, B2 => n1691, C1 => n1171, C2 => 
                           n1688, A => n1017, ZN => n741);
   U2354 : AOI22_X1 port map( A1 => RF_WR_DATAx25x, A2 => n1687, B1 => 
                           RF_RD2_DATA(25), B2 => n1683, ZN => n1017);
   U2355 : OAI221_X1 port map( B1 => n1428, B2 => n1692, C1 => n1184, C2 => 
                           n1689, A => n1041, ZN => n770);
   U2356 : AOI22_X1 port map( A1 => RF_WR_DATAx9x, A2 => n1687, B1 => 
                           RF_RD2_DATA(9), B2 => n1684, ZN => n1041);
   U2357 : OAI221_X1 port map( B1 => n1447, B2 => n1692, C1 => n1166, C2 => 
                           n1689, A => n1030, ZN => n735);
   U2358 : AOI22_X1 port map( A1 => RF_WR_DATAx28x, A2 => n1687, B1 => 
                           RF_RD2_DATA(28), B2 => n1684, ZN => n1030);
   U2359 : OAI221_X1 port map( B1 => n1443, B2 => n1691, C1 => n1172, C2 => 
                           n1688, A => n1020, ZN => n742);
   U2360 : AOI22_X1 port map( A1 => RF_WR_DATAx24x, A2 => n1687, B1 => 
                           RF_RD2_DATA(24), B2 => n1683, ZN => n1020);
   U2361 : OAI221_X1 port map( B1 => n1429, B2 => n1692, C1 => n1186, C2 => 
                           n1689, A => n1055, ZN => n768);
   U2362 : AOI22_X1 port map( A1 => RF_WR_DATAx10x, A2 => n1686, B1 => 
                           RF_RD2_DATA(10), B2 => n1684, ZN => n1055);
   U2363 : OAI221_X1 port map( B1 => n1704, B2 => n1598, C1 => n1419, C2 => 
                           n1701, A => n1068, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_0_port);
   U2364 : AOI22_X1 port map( A1 => RF_WR_DATAx0x, A2 => n1697, B1 => 
                           RF_RD1_DATA(0), B2 => n1694, ZN => n1068);
   U2365 : OAI221_X1 port map( B1 => n1703, B2 => n1587, C1 => n1446, C2 => 
                           n1700, A => n1026, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_27_port);
   U2366 : AOI22_X1 port map( A1 => RF_WR_DATAx27x, A2 => n1698, B1 => 
                           RF_RD1_DATA(27), B2 => n1695, ZN => n1026);
   U2367 : OAI221_X1 port map( B1 => n1703, B2 => n1580, C1 => n1434, C2 => 
                           n1700, A => n1046, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_15_port);
   U2368 : AOI22_X1 port map( A1 => RF_WR_DATAx15x, A2 => n1697, B1 => 
                           RF_RD1_DATA(15), B2 => n1695, ZN => n1046);
   U2369 : OAI221_X1 port map( B1 => n1703, B2 => n1602, C1 => n1433, C2 => 
                           n1700, A => n1043, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_14_port);
   U2370 : AOI22_X1 port map( A1 => RF_WR_DATAx14x, A2 => n1698, B1 => 
                           RF_RD1_DATA(14), B2 => n1695, ZN => n1043);
   U2371 : OAI221_X1 port map( B1 => n1703, B2 => n1605, C1 => n1432, C2 => 
                           n1700, A => n1061, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_13_port);
   U2372 : AOI22_X1 port map( A1 => RF_WR_DATAx13x, A2 => n1697, B1 => 
                           RF_RD1_DATA(13), B2 => n1694, ZN => n1061);
   U2373 : OAI221_X1 port map( B1 => n1703, B2 => n1606, C1 => n1431, C2 => 
                           n1700, A => n1050, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_12_port);
   U2374 : AOI22_X1 port map( A1 => RF_WR_DATAx12x, A2 => n1697, B1 => 
                           RF_RD1_DATA(12), B2 => n1694, ZN => n1050);
   U2375 : OAI221_X1 port map( B1 => n1704, B2 => n1596, C1 => n1424, C2 => 
                           n1701, A => n1074, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_5_port);
   U2376 : AOI22_X1 port map( A1 => RF_WR_DATAx5x, A2 => n1697, B1 => 
                           RF_RD1_DATA(5), B2 => n1694, ZN => n1074);
   U2377 : OAI221_X1 port map( B1 => n1704, B2 => n1581, C1 => n1423, C2 => 
                           n1701, A => n1071, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_4_port);
   U2378 : AOI22_X1 port map( A1 => RF_WR_DATAx4x, A2 => n1697, B1 => 
                           RF_RD1_DATA(4), B2 => n1694, ZN => n1071);
   U2379 : OAI221_X1 port map( B1 => n1702, B2 => n1582, C1 => n1444, C2 => 
                           n1699, A => n1016, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_25_port);
   U2380 : AOI22_X1 port map( A1 => RF_WR_DATAx25x, A2 => n1698, B1 => 
                           RF_RD1_DATA(25), B2 => n1695, ZN => n1016);
   U2381 : NOR2_X1 port map( A1 => n956, A2 => n1244, ZN => n271);
   U2382 : XNOR2_X1 port map( A => n830, B => n831, ZN => n111);
   U2383 : XNOR2_X1 port map( A => n1363, B => n1386, ZN => n830);
   U2384 : OAI21_X1 port map( B1 => n819, B2 => n1659, A => n832, ZN => n831);
   U2385 : OAI21_X1 port map( B1 => n1386, B2 => n1815, A => n1362, ZN => n832)
                           ;
   U2386 : NAND2_X1 port map( A1 => n1241, A2 => n283, ZN => n284);
   U2387 : NAND4_X1 port map( A1 => n1126, A2 => n1127, A3 => n1128, A4 => 
                           n1129, ZN => n1115);
   U2388 : XNOR2_X1 port map( A => n1152, B => n1145, ZN => n1127);
   U2389 : XNOR2_X1 port map( A => n1158, B => n1154, ZN => n1126);
   U2390 : XNOR2_X1 port map( A => n1153, B => n1146, ZN => n1128);
   U2391 : NAND4_X1 port map( A1 => n1102, A2 => n1103, A3 => n1104, A4 => 
                           n1105, ZN => n1093);
   U2392 : XNOR2_X1 port map( A => n1163, B => n1146, ZN => n1102);
   U2393 : XNOR2_X1 port map( A => n1162, B => n1159, ZN => n1104);
   U2394 : XNOR2_X1 port map( A => n1161, B => n1145, ZN => n1103);
   U2395 : XNOR2_X1 port map( A => n836, B => n848, ZN => 
                           DATAPATH_IxSecond_stxjump_target_25_port);
   U2396 : OAI21_X1 port map( B1 => n835, B2 => n1659, A => n849, ZN => n848);
   U2397 : OAI21_X1 port map( B1 => n1386, B2 => n1810, A => n1358, ZN => n849)
                           ;
   U2398 : INV_X1 port map( A => DATAPATH_IxThird_stxALU1xN222, ZN => n1729);
   U2399 : OAI221_X1 port map( B1 => n1702, B2 => n1589, C1 => n1450, C2 => 
                           n1699, A => n1013, ZN => 
                           DATAPATH_IxThird_stxALU1xN222);
   U2400 : AOI22_X1 port map( A1 => RF_WR_DATAx31x, A2 => n1698, B1 => 
                           RF_RD1_DATA(31), B2 => n1695, ZN => n1013);
   U2401 : XNOR2_X1 port map( A => n865, B => n852, ZN => 
                           DATAPATH_IxSecond_stxjump_target_21_port);
   U2402 : OAI21_X1 port map( B1 => n1660, B2 => n181, A => n866, ZN => n865);
   U2403 : OAI21_X1 port map( B1 => n1805, B2 => n1386, A => n1354, ZN => n866)
                           ;
   U2404 : AND2_X1 port map( A1 => n1244, A2 => n956, ZN => n270);
   U2405 : OAI211_X1 port map( C1 => n1405, C2 => n187, A => n188, B => n189, 
                           ZN => n1529);
   U2406 : NAND4_X1 port map( A1 => n1405, A2 => n1632, A3 => n192, A4 => 
                           IRAM_ADD_17_port, ZN => n188);
   U2407 : AOI21_X1 port map( B1 => n1404, B2 => n1632, A => n194, ZN => n187);
   U2408 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_18_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_18_port, ZN 
                           => n189);
   U2409 : INV_X1 port map( A => n1001, ZN => n1903);
   U2410 : OAI221_X1 port map( B1 => n1442, B2 => n1691, C1 => n1174, C2 => 
                           n1688, A => n1002, ZN => n1001);
   U2411 : AOI22_X1 port map( A1 => RF_WR_DATAx23x, A2 => n1687, B1 => 
                           RF_RD2_DATA(23), B2 => n1683, ZN => n1002);
   U2412 : INV_X1 port map( A => n980, ZN => n1908);
   U2413 : OAI221_X1 port map( B1 => n1438, B2 => n1691, C1 => n1177, C2 => 
                           n1688, A => n983, ZN => n980);
   U2414 : AOI22_X1 port map( A1 => RF_WR_DATAx19x, A2 => n1686, B1 => 
                           RF_RD2_DATA(19), B2 => n1683, ZN => n983);
   U2415 : INV_X1 port map( A => n1047, ZN => n1913);
   U2416 : OAI221_X1 port map( B1 => n1434, B2 => n1692, C1 => n1181, C2 => 
                           n1689, A => n1048, ZN => n1047);
   U2417 : AOI22_X1 port map( A1 => RF_WR_DATAx15x, A2 => n1686, B1 => 
                           RF_RD2_DATA(15), B2 => n1684, ZN => n1048);
   U2418 : INV_X1 port map( A => n1058, ZN => n1917);
   U2419 : OAI221_X1 port map( B1 => n1430, B2 => n1692, C1 => n1187, C2 => 
                           n1689, A => n1059, ZN => n1058);
   U2420 : AOI22_X1 port map( A1 => RF_WR_DATAx11x, A2 => n1686, B1 => 
                           RF_RD2_DATA(11), B2 => n1684, ZN => n1059);
   U2421 : INV_X1 port map( A => n1082, ZN => RF_WR_DATAx2x);
   U2422 : OAI22_X1 port map( A1 => n1675, A2 => DATAPATH_IxLMD_DATA_2_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_2_port, ZN 
                           => n1082);
   U2423 : INV_X1 port map( A => n1051, ZN => n1916);
   U2424 : OAI221_X1 port map( B1 => n1431, B2 => n1692, C1 => n1182, C2 => 
                           n1689, A => n1052, ZN => n1051);
   U2425 : AOI22_X1 port map( A1 => RF_WR_DATAx12x, A2 => n1686, B1 => 
                           RF_RD2_DATA(12), B2 => n1684, ZN => n1052);
   U2426 : INV_X1 port map( A => n1070, ZN => RF_WR_DATAx0x);
   U2427 : OAI22_X1 port map( A1 => n1676, A2 => DATAPATH_IxLMD_DATA_0_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_0_port, ZN 
                           => n1070);
   U2428 : INV_X1 port map( A => n1114, ZN => RF_WR_DATAx1x);
   U2429 : OAI22_X1 port map( A1 => n1675, A2 => DATAPATH_IxLMD_DATA_1_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_1_port, ZN 
                           => n1114);
   U2430 : INV_X1 port map( A => n1085, ZN => RF_WR_DATAx3x);
   U2431 : OAI22_X1 port map( A1 => n1675, A2 => DATAPATH_IxLMD_DATA_3_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_3_port, ZN 
                           => n1085);
   U2432 : INV_X1 port map( A => n1073, ZN => RF_WR_DATAx4x);
   U2433 : OAI22_X1 port map( A1 => n1676, A2 => DATAPATH_IxLMD_DATA_4_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_4_port, ZN 
                           => n1073);
   U2434 : INV_X1 port map( A => n1076, ZN => RF_WR_DATAx5x);
   U2435 : OAI22_X1 port map( A1 => n1675, A2 => DATAPATH_IxLMD_DATA_5_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_5_port, ZN 
                           => n1076);
   U2436 : INV_X1 port map( A => n1079, ZN => RF_WR_DATAx6x);
   U2437 : OAI22_X1 port map( A1 => n1675, A2 => DATAPATH_IxLMD_DATA_6_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_6_port, ZN 
                           => n1079);
   U2438 : INV_X1 port map( A => n1067, ZN => RF_WR_DATAx7x);
   U2439 : OAI22_X1 port map( A1 => n1676, A2 => DATAPATH_IxLMD_DATA_7_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_7_port, ZN 
                           => n1067);
   U2440 : INV_X1 port map( A => n1039, ZN => RF_WR_DATAx8x);
   U2441 : OAI22_X1 port map( A1 => n1678, A2 => DATAPATH_IxLMD_DATA_8_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_8_port, ZN 
                           => n1039);
   U2442 : INV_X1 port map( A => n1042, ZN => RF_WR_DATAx9x);
   U2443 : OAI22_X1 port map( A1 => n1677, A2 => DATAPATH_IxLMD_DATA_9_port, B1
                           => n1573, B2 => DATAPATH_IxALUOUT_Data1_9_port, ZN 
                           => n1042);
   U2444 : INV_X1 port map( A => n1056, ZN => RF_WR_DATAx10x);
   U2445 : OAI22_X1 port map( A1 => n1677, A2 => DATAPATH_IxLMD_DATA_10_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_10_port, 
                           ZN => n1056);
   U2446 : INV_X1 port map( A => n1060, ZN => RF_WR_DATAx11x);
   U2447 : OAI22_X1 port map( A1 => n1676, A2 => DATAPATH_IxLMD_DATA_11_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_11_port, 
                           ZN => n1060);
   U2448 : INV_X1 port map( A => n1053, ZN => RF_WR_DATAx12x);
   U2449 : OAI22_X1 port map( A1 => n1677, A2 => DATAPATH_IxLMD_DATA_12_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_12_port, 
                           ZN => n1053);
   U2450 : INV_X1 port map( A => n1063, ZN => RF_WR_DATAx13x);
   U2451 : OAI22_X1 port map( A1 => n1676, A2 => DATAPATH_IxLMD_DATA_13_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_13_port, 
                           ZN => n1063);
   U2452 : INV_X1 port map( A => n1045, ZN => RF_WR_DATAx14x);
   U2453 : OAI22_X1 port map( A1 => n1677, A2 => DATAPATH_IxLMD_DATA_14_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_14_port, 
                           ZN => n1045);
   U2454 : INV_X1 port map( A => n1049, ZN => RF_WR_DATAx15x);
   U2455 : OAI22_X1 port map( A1 => n1677, A2 => DATAPATH_IxLMD_DATA_15_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_15_port, 
                           ZN => n1049);
   U2456 : INV_X1 port map( A => n993, ZN => RF_WR_DATAx16x);
   U2457 : OAI22_X1 port map( A1 => n1680, A2 => DATAPATH_IxLMD_DATA_16_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_16_port, 
                           ZN => n993);
   U2458 : INV_X1 port map( A => n1009, ZN => RF_WR_DATAx17x);
   U2459 : OAI22_X1 port map( A1 => n1679, A2 => DATAPATH_IxLMD_DATA_17_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_17_port, 
                           ZN => n1009);
   U2460 : INV_X1 port map( A => n1006, ZN => RF_WR_DATAx18x);
   U2461 : OAI22_X1 port map( A1 => n1680, A2 => DATAPATH_IxLMD_DATA_18_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_18_port, 
                           ZN => n1006);
   U2462 : INV_X1 port map( A => n986, ZN => RF_WR_DATAx19x);
   U2463 : OAI22_X1 port map( A1 => n1681, A2 => DATAPATH_IxLMD_DATA_19_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_19_port, 
                           ZN => n986);
   U2464 : INV_X1 port map( A => n996, ZN => RF_WR_DATAx20x);
   U2465 : OAI22_X1 port map( A1 => n1680, A2 => DATAPATH_IxLMD_DATA_20_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_20_port, 
                           ZN => n996);
   U2466 : INV_X1 port map( A => n999, ZN => RF_WR_DATAx21x);
   U2467 : OAI22_X1 port map( A1 => n1680, A2 => DATAPATH_IxLMD_DATA_21_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_21_port, 
                           ZN => n999);
   U2468 : INV_X1 port map( A => n990, ZN => RF_WR_DATAx22x);
   U2469 : OAI22_X1 port map( A1 => n1681, A2 => DATAPATH_IxLMD_DATA_22_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_22_port, 
                           ZN => n990);
   U2470 : INV_X1 port map( A => n1003, ZN => RF_WR_DATAx23x);
   U2471 : OAI22_X1 port map( A1 => n1680, A2 => DATAPATH_IxLMD_DATA_23_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_23_port, 
                           ZN => n1003);
   U2472 : INV_X1 port map( A => n1021, ZN => RF_WR_DATAx24x);
   U2473 : OAI22_X1 port map( A1 => n1679, A2 => DATAPATH_IxLMD_DATA_24_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_24_port, 
                           ZN => n1021);
   U2474 : INV_X1 port map( A => n1018, ZN => RF_WR_DATAx25x);
   U2475 : OAI22_X1 port map( A1 => n1679, A2 => DATAPATH_IxLMD_DATA_25_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_25_port, 
                           ZN => n1018);
   U2476 : INV_X1 port map( A => n1025, ZN => RF_WR_DATAx26x);
   U2477 : OAI22_X1 port map( A1 => n1678, A2 => DATAPATH_IxLMD_DATA_26_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_26_port, 
                           ZN => n1025);
   U2478 : INV_X1 port map( A => n1028, ZN => RF_WR_DATAx27x);
   U2479 : OAI22_X1 port map( A1 => n1678, A2 => DATAPATH_IxLMD_DATA_27_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_27_port, 
                           ZN => n1028);
   U2480 : INV_X1 port map( A => n1031, ZN => RF_WR_DATAx28x);
   U2481 : OAI22_X1 port map( A1 => n1678, A2 => DATAPATH_IxLMD_DATA_28_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_28_port, 
                           ZN => n1031);
   U2482 : INV_X1 port map( A => n1012, ZN => RF_WR_DATAx30x);
   U2483 : OAI22_X1 port map( A1 => n1679, A2 => DATAPATH_IxLMD_DATA_30_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_30_port, 
                           ZN => n1012);
   U2484 : INV_X1 port map( A => n1015, ZN => RF_WR_DATAx31x);
   U2485 : OAI22_X1 port map( A1 => n1679, A2 => DATAPATH_IxLMD_DATA_31_port, 
                           B1 => n1674, B2 => DATAPATH_IxALUOUT_Data1_31_port, 
                           ZN => n1015);
   U2486 : INV_X1 port map( A => n1034, ZN => RF_WR_DATAx29x);
   U2487 : OAI22_X1 port map( A1 => n1678, A2 => DATAPATH_IxLMD_DATA_29_port, 
                           B1 => n1573, B2 => DATAPATH_IxALUOUT_Data1_29_port, 
                           ZN => n1034);
   U2488 : INV_X1 port map( A => n945, ZN => n1833);
   U2489 : AOI22_X1 port map( A1 => n897, A2 => n1366, B1 => n1847, B2 => n1376
                           , ZN => n945);
   U2490 : AND4_X1 port map( A1 => n1155, A2 => n1156, A3 => n1154, A4 => n1132
                           , ZN => n1120);
   U2491 : AND2_X1 port map( A1 => n1153, A2 => n1152, ZN => n1132);
   U2492 : AND4_X1 port map( A1 => n1164, A2 => n1165, A3 => n1163, A4 => n1108
                           , ZN => n1096);
   U2493 : AND2_X1 port map( A1 => n1162, A2 => n1161, ZN => n1108);
   U2494 : OAI221_X1 port map( B1 => n1647, B2 => n1816, C1 => n1226, C2 => 
                           n1649, A => n174, ZN => n1527);
   U2495 : AOI21_X1 port map( B1 => n175, B2 => IRAM_ADD_20_port, A => n177, ZN
                           => n174);
   U2496 : INV_X1 port map( A => n1292, ZN => n1816);
   U2497 : OAI21_X1 port map( B1 => n1646, B2 => IRAM_ADD_19_port, A => n179, 
                           ZN => n175);
   U2498 : OAI221_X1 port map( B1 => n1237, B2 => n1650, C1 => n1812, C2 => 
                           n1648, A => n96, ZN => n1516);
   U2499 : AOI21_X1 port map( B1 => n97, B2 => IRAM_ADD_31_port, A => n99, ZN 
                           => n96);
   U2500 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_31_port, ZN 
                           => n1812);
   U2501 : OAI21_X1 port map( B1 => n1645, B2 => IRAM_ADD_30_port, A => n103, 
                           ZN => n97);
   U2502 : OAI221_X1 port map( B1 => n1236, B2 => n1649, C1 => n1813, C2 => 
                           n1647, A => n105, ZN => n1517);
   U2503 : AOI22_X1 port map( A1 => n106, A2 => n1417, B1 => n1764, B2 => 
                           IRAM_ADD_30_port, ZN => n105);
   U2504 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_30_port, ZN 
                           => n1813);
   U2505 : INV_X1 port map( A => n103, ZN => n1764);
   U2506 : INV_X1 port map( A => n292, ZN => n1854);
   U2507 : AOI211_X1 port map( C1 => n1830, C2 => n1372, A => n896, B => n1350,
                           ZN => n878);
   U2508 : AOI211_X1 port map( C1 => n1847, C2 => n1210, A => n882, B => n1622,
                           ZN => n916);
   U2509 : AOI211_X1 port map( C1 => n1830, C2 => n1374, A => n896, B => n1352,
                           ZN => n872);
   U2510 : AOI21_X1 port map( B1 => n1632, B2 => n1414, A => n124, ZN => n119);
   U2511 : NOR4_X1 port map( A1 => n1417, A2 => n1645, A3 => n101, A4 => 
                           IRAM_ADD_31_port, ZN => n99);
   U2512 : NOR4_X1 port map( A1 => n1412, A2 => n132, A3 => n1644, A4 => 
                           IRAM_ADD_26_port, ZN => n137);
   U2513 : NOR4_X1 port map( A1 => n1406, A2 => n172, A3 => n1644, A4 => 
                           IRAM_ADD_20_port, ZN => n177);
   U2514 : NOR4_X1 port map( A1 => n1402, A2 => n198, A3 => n1644, A4 => 
                           IRAM_ADD_16_port, ZN => n203);
   U2515 : AOI21_X1 port map( B1 => n1632, B2 => n1390, A => n267, ZN => n266);
   U2516 : OAI222_X1 port map( A1 => n1213, A2 => n1650, B1 => n1387, B2 => 
                           n285, C1 => n1338, C2 => n1648, ZN => n1547);
   U2517 : OAI222_X1 port map( A1 => n1648, A2 => n49, B1 => n1388, B2 => n285,
                           C1 => n1214, C2 => n1650, ZN => n1546);
   U2518 : OAI21_X1 port map( B1 => n291, B2 => n1211, A => n292, ZN => n165);
   U2519 : OAI211_X1 port map( C1 => n1372, C2 => n897, A => n1830, B => n1350,
                           ZN => n877);
   U2520 : NOR2_X1 port map( A1 => n1197, A2 => n1298, ZN => n298);
   U2521 : AOI21_X1 port map( B1 => RF_RD1_ADD_4_port, B2 => n1847, A => n882, 
                           ZN => n867);
   U2522 : OAI221_X1 port map( B1 => n1222, B2 => n1650, C1 => n1648, C2 => 
                           n206, A => n207, ZN => n1532);
   U2523 : AOI21_X1 port map( B1 => n1760, B2 => IRAM_ADD_15_port, A => n209, 
                           ZN => n207);
   U2524 : INV_X1 port map( A => n205, ZN => n1760);
   U2525 : NOR3_X1 port map( A1 => IRAM_ADD_15_port, A2 => n198, A3 => n1645, 
                           ZN => n209);
   U2526 : OAI221_X1 port map( B1 => n1221, B2 => n1650, C1 => n217, C2 => 
                           n1648, A => n218, ZN => n1534);
   U2527 : AOI21_X1 port map( B1 => n216, B2 => IRAM_ADD_13_port, A => n219, ZN
                           => n218);
   U2528 : NOR3_X1 port map( A1 => IRAM_ADD_13_port, A2 => n1973, A3 => n1645, 
                           ZN => n219);
   U2529 : OAI221_X1 port map( B1 => n1220, B2 => n1650, C1 => n1832, C2 => 
                           n1648, A => n228, ZN => n1536);
   U2530 : AOI21_X1 port map( B1 => n226, B2 => IRAM_ADD_11_port, A => n229, ZN
                           => n228);
   U2531 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_11_port, ZN 
                           => n1832);
   U2532 : NOR3_X1 port map( A1 => IRAM_ADD_11_port, A2 => n1974, A3 => n1645, 
                           ZN => n229);
   U2533 : OAI221_X1 port map( B1 => n1219, B2 => n1650, C1 => n1648, C2 => 
                           n237, A => n238, ZN => n1538);
   U2534 : AOI21_X1 port map( B1 => n236, B2 => IRAM_ADD_9_port, A => n239, ZN 
                           => n238);
   U2535 : NOR3_X1 port map( A1 => IRAM_ADD_9_port, A2 => n1975, A3 => n1645, 
                           ZN => n239);
   U2536 : OAI221_X1 port map( B1 => n1218, B2 => n1650, C1 => n1834, C2 => 
                           n1648, A => n250, ZN => n1540);
   U2537 : AOI21_X1 port map( B1 => n248, B2 => IRAM_ADD_7_port, A => n251, ZN 
                           => n250);
   U2538 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_7_port, ZN =>
                           n1834);
   U2539 : NOR3_X1 port map( A1 => IRAM_ADD_7_port, A2 => n1976, A3 => n1645, 
                           ZN => n251);
   U2540 : OAI221_X1 port map( B1 => n1217, B2 => n1650, C1 => n1835, C2 => 
                           n1648, A => n260, ZN => n1542);
   U2541 : AOI21_X1 port map( B1 => n258, B2 => IRAM_ADD_5_port, A => n261, ZN 
                           => n260);
   U2542 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_5_port, ZN =>
                           n1835);
   U2543 : NOR3_X1 port map( A1 => IRAM_ADD_5_port, A2 => n1977, A3 => n1644, 
                           ZN => n261);
   U2544 : OAI221_X1 port map( B1 => n1215, B2 => n1650, C1 => n1840, C2 => 
                           n1648, A => n273, ZN => n1544);
   U2545 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_3_port, ZN =>
                           n1840);
   U2546 : AOI21_X1 port map( B1 => n267, B2 => IRAM_ADD_3_port, A => n275, ZN 
                           => n273);
   U2547 : NOR3_X1 port map( A1 => IRAM_ADD_3_port, A2 => n1389, A3 => n1644, 
                           ZN => n275);
   U2548 : OAI221_X1 port map( B1 => n1644, B2 => IRAM_ADD_2_port, C1 => n1648,
                           C2 => n1842, A => n278, ZN => n1545);
   U2549 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_2_port, B1 => n109, 
                           B2 => IRAM_ADD_2_port, ZN => n278);
   U2550 : INV_X1 port map( A => n1296, ZN => n1842);
   U2551 : OAI211_X1 port map( C1 => n1373, C2 => n897, A => n1830, B => n1351,
                           ZN => n894);
   U2552 : OAI21_X1 port map( B1 => n294, B2 => n1924, A => n1793, ZN => n296);
   U2553 : INV_X1 port map( A => CU_Ixcw_LUT_16_port, ZN => n1793);
   U2554 : OAI21_X1 port map( B1 => n1924, B2 => n294, A => n1212, ZN => n292);
   U2555 : OAI211_X1 port map( C1 => n1374, C2 => n897, A => n1830, B => n1352,
                           ZN => n887);
   U2556 : OAI22_X1 port map( A1 => n1727, A2 => n1575, B1 => n1362, B2 => 
                           n1721, ZN => n1458);
   U2557 : OAI22_X1 port map( A1 => n1726, A2 => n1576, B1 => n1358, B2 => 
                           n1721, ZN => n1466);
   U2558 : OAI22_X1 port map( A1 => n1726, A2 => n1577, B1 => n1354, B2 => 
                           n1721, ZN => n1474);
   U2559 : OAI22_X1 port map( A1 => n1723, A2 => n1592, B1 => n1343, B2 => 
                           n1720, ZN => n1498);
   U2560 : OAI22_X1 port map( A1 => n1723, A2 => n1594, B1 => n1344, B2 => 
                           n1720, ZN => n1496);
   U2561 : OAI22_X1 port map( A1 => n1727, A2 => n1574, B1 => n1363, B2 => 
                           n1721, ZN => n1456);
   U2562 : OAI22_X1 port map( A1 => n1727, A2 => n1582, B1 => n1359, B2 => 
                           n1720, ZN => n1464);
   U2563 : OAI22_X1 port map( A1 => n1726, A2 => n1583, B1 => n1355, B2 => 
                           n1721, ZN => n1472);
   U2564 : XNOR2_X1 port map( A => n867, B => n1353, ZN => n869);
   U2565 : OAI22_X1 port map( A1 => n1723, A2 => n1595, B1 => n1342, B2 => 
                           n1721, ZN => n1502);
   U2566 : OAI22_X1 port map( A1 => n1723, A2 => n1596, B1 => n1341, B2 => 
                           n1721, ZN => n1504);
   U2567 : OAI22_X1 port map( A1 => n1722, A2 => n1597, B1 => n1340, B2 => 
                           n1721, ZN => n1508);
   U2568 : OAI22_X1 port map( A1 => n1722, A2 => n1598, B1 => n1338, B2 => 
                           n1721, ZN => n1514);
   U2569 : OAI22_X1 port map( A1 => n1722, A2 => n1599, B1 => n1339, B2 => 
                           n1721, ZN => n1512);
   U2570 : OAI22_X1 port map( A1 => n1725, A2 => n1600, B1 => n1353, B2 => 
                           n1720, ZN => n1476);
   U2571 : OAI22_X1 port map( A1 => n1724, A2 => n1601, B1 => n1346, B2 => 
                           n1720, ZN => n1492);
   U2572 : OAI22_X1 port map( A1 => n1728, A2 => n1584, B1 => n1364, B2 => 
                           n1720, ZN => n1454);
   U2573 : OAI22_X1 port map( A1 => n1727, A2 => n1585, B1 => n1360, B2 => 
                           n1721, ZN => n1462);
   U2574 : OAI22_X1 port map( A1 => n1726, A2 => n1586, B1 => n1356, B2 => 
                           n1720, ZN => n1470);
   U2575 : OAI22_X1 port map( A1 => n1727, A2 => n1587, B1 => n1361, B2 => 
                           n1721, ZN => n1460);
   U2576 : OAI22_X1 port map( A1 => n1726, A2 => n1588, B1 => n1357, B2 => 
                           n1720, ZN => n1468);
   U2577 : OAI22_X1 port map( A1 => n1724, A2 => n1602, B1 => n1349, B2 => 
                           n1720, ZN => n1486);
   U2578 : OAI22_X1 port map( A1 => n1725, A2 => n1603, B1 => n1352, B2 => 
                           n1720, ZN => n1478);
   U2579 : OAI22_X1 port map( A1 => n1725, A2 => n1604, B1 => n1351, B2 => 
                           n1720, ZN => n1480);
   U2580 : OAI22_X1 port map( A1 => n1725, A2 => n1593, B1 => n1350, B2 => 
                           n1720, ZN => n1482);
   U2581 : OAI22_X1 port map( A1 => n1724, A2 => n1605, B1 => n1348, B2 => 
                           n1720, ZN => n1488);
   U2582 : OAI22_X1 port map( A1 => n1724, A2 => n1606, B1 => n1347, B2 => 
                           n1720, ZN => n1490);
   U2583 : OAI22_X1 port map( A1 => n1724, A2 => n1607, B1 => n1345, B2 => 
                           n1720, ZN => n1494);
   U2584 : OAI22_X1 port map( A1 => n1728, A2 => n1589, B1 => n1365, B2 => 
                           n1721, ZN => n1452);
   U2585 : AOI22_X1 port map( A1 => n1837, A2 => n1963, B1 => n1384, B2 => 
                           n1343, ZN => n792);
   U2586 : INV_X1 port map( A => n794, ZN => n1963);
   U2587 : INV_X1 port map( A => n899, ZN => n1826);
   U2588 : AOI211_X1 port map( C1 => n1830, C2 => n1373, A => n896, B => n1351,
                           ZN => n899);
   U2589 : OAI211_X1 port map( C1 => n1401, C2 => n211, A => n212, B => n213, 
                           ZN => n1533);
   U2590 : NAND4_X1 port map( A1 => n1401, A2 => n1632, A3 => n214, A4 => 
                           IRAM_ADD_13_port, ZN => n212);
   U2591 : AOI21_X1 port map( B1 => n1400, B2 => n1632, A => n216, ZN => n211);
   U2592 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_14_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_14_port, ZN 
                           => n213);
   U2593 : OAI211_X1 port map( C1 => n1399, C2 => n221, A => n222, B => n223, 
                           ZN => n1535);
   U2594 : NAND4_X1 port map( A1 => n1399, A2 => n1632, A3 => n224, A4 => 
                           IRAM_ADD_11_port, ZN => n222);
   U2595 : AOI21_X1 port map( B1 => n1398, B2 => n1632, A => n226, ZN => n221);
   U2596 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_12_port, B1 => 
                           DATAPATH_IxSecond_stxjump_target_12_port, B2 => n191
                           , ZN => n223);
   U2597 : OAI211_X1 port map( C1 => n1397, C2 => n231, A => n232, B => n233, 
                           ZN => n1537);
   U2598 : NAND4_X1 port map( A1 => n1397, A2 => n1632, A3 => n234, A4 => 
                           IRAM_ADD_9_port, ZN => n232);
   U2599 : AOI21_X1 port map( B1 => n1396, B2 => n1632, A => n236, ZN => n231);
   U2600 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_10_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_10_port, ZN 
                           => n233);
   U2601 : OAI211_X1 port map( C1 => n1395, C2 => n241, A => n242, B => n243, 
                           ZN => n1539);
   U2602 : NAND4_X1 port map( A1 => n1395, A2 => n1632, A3 => n246, A4 => 
                           IRAM_ADD_7_port, ZN => n242);
   U2603 : AOI21_X1 port map( B1 => n1394, B2 => n1632, A => n248, ZN => n241);
   U2604 : AOI22_X1 port map( A1 => n1291, A2 => n191, B1 => n190, B2 => 
                           DATAPATH_IxSecond_stxBR_target_8_port, ZN => n243);
   U2605 : OAI211_X1 port map( C1 => n1393, C2 => n253, A => n254, B => n255, 
                           ZN => n1541);
   U2606 : NAND4_X1 port map( A1 => n1393, A2 => n1632, A3 => n256, A4 => 
                           IRAM_ADD_5_port, ZN => n254);
   U2607 : AOI21_X1 port map( B1 => n1392, B2 => n1632, A => n258, ZN => n253);
   U2608 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_6_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_6_port, ZN =>
                           n255);
   U2609 : NOR2_X1 port map( A1 => n1207, A2 => n291, ZN => RF_RD2_EN);
   U2610 : NOR2_X1 port map( A1 => n1206, A2 => n291, ZN => RF_RD1_EN);
   U2611 : OAI21_X1 port map( B1 => n1371, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_15_port);
   U2612 : OAI21_X1 port map( B1 => n1372, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_16_port);
   U2613 : OAI21_X1 port map( B1 => n1373, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_17_port);
   U2614 : OAI21_X1 port map( B1 => n1374, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_18_port);
   U2615 : OAI21_X1 port map( B1 => n1375, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_19_port);
   U2616 : OAI21_X1 port map( B1 => n1376, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_20_port);
   U2617 : OAI21_X1 port map( B1 => n1377, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_21_port);
   U2618 : OAI21_X1 port map( B1 => n1378, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_22_port);
   U2619 : OAI21_X1 port map( B1 => n1379, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_23_port);
   U2620 : OAI21_X1 port map( B1 => n1380, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_24_port);
   U2621 : OAI21_X1 port map( B1 => n1381, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_25_port);
   U2622 : OAI21_X1 port map( B1 => n1382, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_26_port);
   U2623 : OAI21_X1 port map( B1 => n1383, B2 => n1640, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_27_port);
   U2624 : OAI21_X1 port map( B1 => n1384, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_28_port);
   U2625 : OAI21_X1 port map( B1 => n1385, B2 => n963, A => n1848, ZN => 
                           DATAPATH_IxSecond_stximm_extended_30_port);
   U2626 : OR3_X1 port map( A1 => n291, A2 => n1205, A3 => n1849, ZN => n962);
   U2627 : NAND2_X1 port map( A1 => CU_Ixcw2_i_10_port, A2 => n1850, ZN => 
                           n1451);
   U2628 : BUF_X1 port map( A => n1337, Z => n1661);
   U2629 : OAI221_X1 port map( B1 => n1647, B2 => n48, C1 => n1216, C2 => n1649
                           , A => n262, ZN => n1543);
   U2630 : AOI21_X1 port map( B1 => n1759, B2 => IRAM_ADD_4_port, A => n265, ZN
                           => n262);
   U2631 : NOR4_X1 port map( A1 => n1389, A2 => n1390, A3 => n1644, A4 => 
                           IRAM_ADD_4_port, ZN => n265);
   U2632 : INV_X1 port map( A => n266, ZN => n1759);
   U2633 : AOI21_X1 port map( B1 => n279, B2 => n280, A => n1843, ZN => n1296);
   U2634 : OAI21_X1 port map( B1 => n283, B2 => n1241, A => n284, ZN => n280);
   U2635 : INV_X1 port map( A => n282, ZN => n1843);
   U2636 : AND2_X1 port map( A1 => CU_Ixcw2_i_11_port, A2 => n1850, ZN => n1635
                           );
   U2637 : OAI21_X1 port map( B1 => n1205, B2 => n291, A => n1451, ZN => n961);
   U2638 : NOR3_X1 port map( A1 => n1800, A2 => IRAM_DOUT(3), A3 => n1799, ZN 
                           => n1137);
   U2639 : NOR3_X1 port map( A1 => n1390, A2 => n1389, A3 => n1391, ZN => n256)
                           ;
   U2640 : NOR3_X1 port map( A1 => n1403, A2 => n1402, A3 => n198, ZN => n192);
   U2641 : NOR3_X1 port map( A1 => n1399, A2 => n1398, A3 => n1974, ZN => n214)
                           ;
   U2642 : NOR3_X1 port map( A1 => n1397, A2 => n1396, A3 => n1975, ZN => n224)
                           ;
   U2643 : NOR3_X1 port map( A1 => n1395, A2 => n1394, A3 => n1976, ZN => n234)
                           ;
   U2644 : NOR3_X1 port map( A1 => n1393, A2 => n1392, A3 => n1977, ZN => n246)
                           ;
   U2645 : NAND2_X1 port map( A1 => n1205, A2 => n1849, ZN => n963);
   U2646 : NAND2_X1 port map( A1 => n1205, A2 => n1849, ZN => n1640);
   U2647 : NOR3_X1 port map( A1 => n1413, A2 => n1412, A3 => n132, ZN => n118);
   U2648 : NAND4_X1 port map( A1 => IRAM_DOUT(2), A2 => IRAM_DOUT(6), A3 => 
                           IRAM_DOUT(3), A4 => n1141, ZN => n1134);
   U2649 : NOR4_X1 port map( A1 => IRAM_DOUT(4), A2 => n1800, A3 => n1799, A4 
                           => n1796, ZN => n1141);
   U2650 : OR3_X1 port map( A1 => IRAM_DOUT(2), A2 => IRAM_DOUT(5), A3 => n1794
                           , ZN => n1139);
   U2651 : OAI21_X1 port map( B1 => n1140, B2 => n1794, A => n1134, ZN => 
                           CU_IxN23);
   U2652 : AOI22_X1 port map( A1 => n27, A2 => n1797, B1 => IRAM_DOUT(4), B2 =>
                           n1796, ZN => n1140);
   U2653 : NOR2_X1 port map( A1 => n1796, A2 => IRAM_DOUT(2), ZN => n27);
   U2654 : NOR3_X1 port map( A1 => n1407, A2 => n1406, A3 => n172, ZN => n171);
   U2655 : NOR2_X1 port map( A1 => n1343, A2 => n1384, ZN => n794);
   U2656 : NOR2_X1 port map( A1 => n1385, A2 => n1345, ZN => n933);
   U2657 : NOR2_X1 port map( A1 => n1341, A2 => n1381, ZN => n811);
   U2658 : NAND4_X1 port map( A1 => IRAM_DOUT(6), A2 => n27, A3 => n1137, A4 =>
                           n1797, ZN => n26);
   U2659 : NOR2_X1 port map( A1 => n1408, A2 => n1971, ZN => n164);
   U2660 : XNOR2_X1 port map( A => n1344, B => n1624, ZN => n791);
   U2661 : OAI22_X1 port map( A1 => n1643, A2 => n1610, B1 => n1389, B2 => 
                           n1719, ZN => n1511);
   U2662 : OAI22_X1 port map( A1 => n1355, A2 => n1642, B1 => n1408, B2 => 
                           n1717, ZN => n1473);
   U2663 : OAI22_X1 port map( A1 => n1340, A2 => n1641, B1 => n1390, B2 => 
                           n1719, ZN => n1509);
   U2664 : OAI22_X1 port map( A1 => n1346, A2 => n1641, B1 => n1398, B2 => 
                           n1718, ZN => n1493);
   U2665 : OAI22_X1 port map( A1 => n1344, A2 => n1641, B1 => n1396, B2 => 
                           n1718, ZN => n1497);
   U2666 : OAI22_X1 port map( A1 => n1643, A2 => n1611, B1 => n1394, B2 => 
                           n1719, ZN => n1501);
   U2667 : OAI22_X1 port map( A1 => n1341, A2 => n1641, B1 => n1392, B2 => 
                           n1719, ZN => n1505);
   U2668 : OAI22_X1 port map( A1 => n1351, A2 => n1642, B1 => n1404, B2 => 
                           n1718, ZN => n1481);
   U2669 : OAI22_X1 port map( A1 => n1348, A2 => n1641, B1 => n1400, B2 => 
                           n1718, ZN => n1489);
   U2670 : OAI22_X1 port map( A1 => n1359, A2 => n1642, B1 => n1412, B2 => 
                           n1717, ZN => n1465);
   U2671 : OAI22_X1 port map( A1 => n1353, A2 => n1642, B1 => n1406, B2 => 
                           n1718, ZN => n1477);
   U2672 : OAI22_X1 port map( A1 => n1643, A2 => n1616, B1 => n1402, B2 => 
                           n1718, ZN => n1485);
   U2673 : OAI22_X1 port map( A1 => n1357, A2 => n1642, B1 => n1410, B2 => 
                           n1717, ZN => n1469);
   U2674 : OAI22_X1 port map( A1 => n1364, A2 => n1643, B1 => n1417, B2 => 
                           n1717, ZN => n1455);
   U2675 : OAI22_X1 port map( A1 => n1361, A2 => n1643, B1 => n1414, B2 => 
                           n1717, ZN => n1461);
   U2676 : OAI22_X1 port map( A1 => n1347, A2 => n1641, B1 => n1399, B2 => 
                           n1718, ZN => n1491);
   U2677 : OAI22_X1 port map( A1 => n1345, A2 => n1641, B1 => n1397, B2 => 
                           n1718, ZN => n1495);
   U2678 : OAI22_X1 port map( A1 => n1343, A2 => n1641, B1 => n1395, B2 => 
                           n1718, ZN => n1499);
   U2679 : OAI22_X1 port map( A1 => n1342, A2 => n1641, B1 => n1393, B2 => 
                           n1719, ZN => n1503);
   U2680 : OAI22_X1 port map( A1 => n1352, A2 => n1642, B1 => n1405, B2 => 
                           n1718, ZN => n1479);
   U2681 : OAI22_X1 port map( A1 => n1349, A2 => n1641, B1 => n1401, B2 => 
                           n1718, ZN => n1487);
   U2682 : OAI22_X1 port map( A1 => n1356, A2 => n1642, B1 => n1409, B2 => 
                           n1717, ZN => n1471);
   U2683 : OAI22_X1 port map( A1 => n1643, A2 => n1620, B1 => n1391, B2 => 
                           n1719, ZN => n1507);
   U2684 : OAI22_X1 port map( A1 => n1338, A2 => n1641, B1 => n1387, B2 => 
                           n1719, ZN => n1515);
   U2685 : OAI22_X1 port map( A1 => n1339, A2 => n1641, B1 => n1388, B2 => 
                           n1719, ZN => n1513);
   U2686 : OAI22_X1 port map( A1 => n1376, A2 => n961, B1 => n1366, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_0_port);
   U2687 : OAI22_X1 port map( A1 => n1377, A2 => n961, B1 => n1367, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_1_port);
   U2688 : OAI22_X1 port map( A1 => n1378, A2 => n961, B1 => n1368, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_2_port);
   U2689 : OAI22_X1 port map( A1 => n1379, A2 => n961, B1 => n1369, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_3_port);
   U2690 : OAI22_X1 port map( A1 => n1360, A2 => n1642, B1 => n1413, B2 => 
                           n1717, ZN => n1463);
   U2691 : OAI22_X1 port map( A1 => n1354, A2 => n1642, B1 => n1407, B2 => 
                           n1717, ZN => n1475);
   U2692 : OAI22_X1 port map( A1 => n1350, A2 => n1642, B1 => n1403, B2 => 
                           n1718, ZN => n1483);
   U2693 : OAI22_X1 port map( A1 => n1358, A2 => n1642, B1 => n1411, B2 => 
                           n1717, ZN => n1467);
   U2694 : OAI22_X1 port map( A1 => n1380, A2 => n961, B1 => n1370, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_4_port);
   U2695 : OAI22_X1 port map( A1 => n1363, A2 => n1643, B1 => n1416, B2 => 
                           n1717, ZN => n1457);
   U2696 : NOR2_X1 port map( A1 => n1382, A2 => n1342, ZN => n805);
   U2697 : OAI22_X1 port map( A1 => n1366, A2 => n1714, B1 => n1712, B2 => 
                           n1792, ZN => n1572);
   U2698 : INV_X1 port map( A => IRAM_DOUT(7), ZN => n1792);
   U2699 : OAI22_X1 port map( A1 => n1367, A2 => n1714, B1 => n1713, B2 => 
                           n1791, ZN => n1571);
   U2700 : INV_X1 port map( A => IRAM_DOUT(8), ZN => n1791);
   U2701 : OAI22_X1 port map( A1 => n1368, A2 => n1714, B1 => n1713, B2 => 
                           n1790, ZN => n1570);
   U2702 : INV_X1 port map( A => IRAM_DOUT(9), ZN => n1790);
   U2703 : OAI22_X1 port map( A1 => n1369, A2 => n1714, B1 => n1713, B2 => 
                           n1789, ZN => n1569);
   U2704 : INV_X1 port map( A => IRAM_DOUT(10), ZN => n1789);
   U2705 : OAI22_X1 port map( A1 => n1370, A2 => n1714, B1 => n1713, B2 => 
                           n1788, ZN => n1568);
   U2706 : INV_X1 port map( A => IRAM_DOUT(11), ZN => n1788);
   U2707 : OAI22_X1 port map( A1 => n1371, A2 => n1714, B1 => n1713, B2 => 
                           n1784, ZN => n1564);
   U2708 : INV_X1 port map( A => IRAM_DOUT(15), ZN => n1784);
   U2709 : OAI22_X1 port map( A1 => n1372, A2 => n1714, B1 => n1713, B2 => 
                           n1783, ZN => n1563);
   U2710 : INV_X1 port map( A => IRAM_DOUT(16), ZN => n1783);
   U2711 : OAI22_X1 port map( A1 => n1373, A2 => n1714, B1 => n1713, B2 => 
                           n1782, ZN => n1562);
   U2712 : INV_X1 port map( A => IRAM_DOUT(17), ZN => n1782);
   U2713 : OAI22_X1 port map( A1 => n1374, A2 => n1715, B1 => n1713, B2 => 
                           n1781, ZN => n1561);
   U2714 : INV_X1 port map( A => IRAM_DOUT(18), ZN => n1781);
   U2715 : OAI22_X1 port map( A1 => n1375, A2 => n1715, B1 => n1713, B2 => 
                           n1780, ZN => n1560);
   U2716 : INV_X1 port map( A => IRAM_DOUT(19), ZN => n1780);
   U2717 : OAI22_X1 port map( A1 => n1376, A2 => n1715, B1 => n1713, B2 => 
                           n1779, ZN => n1559);
   U2718 : INV_X1 port map( A => IRAM_DOUT(20), ZN => n1779);
   U2719 : OAI22_X1 port map( A1 => n1377, A2 => n1715, B1 => n1713, B2 => 
                           n1778, ZN => n1558);
   U2720 : INV_X1 port map( A => IRAM_DOUT(21), ZN => n1778);
   U2721 : OAI22_X1 port map( A1 => n1378, A2 => n1715, B1 => n1713, B2 => 
                           n1777, ZN => n1557);
   U2722 : INV_X1 port map( A => IRAM_DOUT(22), ZN => n1777);
   U2723 : OAI22_X1 port map( A1 => n1379, A2 => n1715, B1 => n1712, B2 => 
                           n1776, ZN => n1556);
   U2724 : INV_X1 port map( A => IRAM_DOUT(23), ZN => n1776);
   U2725 : OAI22_X1 port map( A1 => n1380, A2 => n1715, B1 => n1712, B2 => 
                           n1775, ZN => n1555);
   U2726 : INV_X1 port map( A => IRAM_DOUT(24), ZN => n1775);
   U2727 : OAI22_X1 port map( A1 => n1381, A2 => n1715, B1 => n1712, B2 => 
                           n1774, ZN => n1554);
   U2728 : INV_X1 port map( A => IRAM_DOUT(25), ZN => n1774);
   U2729 : OAI22_X1 port map( A1 => n1382, A2 => n1715, B1 => n1712, B2 => 
                           n1773, ZN => n1553);
   U2730 : INV_X1 port map( A => IRAM_DOUT(26), ZN => n1773);
   U2731 : OAI22_X1 port map( A1 => n1383, A2 => n1715, B1 => n1712, B2 => 
                           n1772, ZN => n1552);
   U2732 : INV_X1 port map( A => IRAM_DOUT(27), ZN => n1772);
   U2733 : OAI22_X1 port map( A1 => n1384, A2 => n1715, B1 => n1712, B2 => 
                           n1771, ZN => n1551);
   U2734 : INV_X1 port map( A => IRAM_DOUT(28), ZN => n1771);
   U2735 : OAI22_X1 port map( A1 => n1624, A2 => n1715, B1 => n1712, B2 => 
                           n1770, ZN => n1550);
   U2736 : INV_X1 port map( A => IRAM_DOUT(29), ZN => n1770);
   U2737 : OAI22_X1 port map( A1 => n1385, A2 => n1716, B1 => n1712, B2 => 
                           n1769, ZN => n1549);
   U2738 : INV_X1 port map( A => IRAM_DOUT(30), ZN => n1769);
   U2739 : OAI22_X1 port map( A1 => n1386, A2 => n1716, B1 => n1713, B2 => 
                           n1768, ZN => n1548);
   U2740 : INV_X1 port map( A => IRAM_DOUT(31), ZN => n1768);
   U2741 : OAI22_X1 port map( A1 => n1365, A2 => n1642, B1 => n1418, B2 => 
                           n1717, ZN => n1453);
   U2742 : OAI22_X1 port map( A1 => n1362, A2 => n1643, B1 => n1415, B2 => 
                           n1717, ZN => n1459);
   U2743 : NOR2_X1 port map( A1 => n1624, A2 => n1344, ZN => n949);
   U2744 : NOR2_X1 port map( A1 => n1798, A2 => IRAM_DOUT(6), ZN => n1138);
   U2745 : INV_X1 port map( A => n1137, ZN => n1798);
   U2746 : INV_X1 port map( A => IRAM_DOUT(4), ZN => n1797);
   U2747 : INV_X1 port map( A => IRAM_DOUT(5), ZN => n1796);
   U2748 : NAND2_X1 port map( A1 => n1341, A2 => n1381, ZN => n809);
   U2749 : AND2_X1 port map( A1 => n1345, A2 => n1385, ZN => n941);
   U2750 : OR2_X1 port map( A1 => n110, A2 => n1416, ZN => n101);
   U2751 : NOR2_X1 port map( A1 => n1198, A2 => n291, ZN => CU_Ixcw2_0_port);
   U2752 : NOR2_X1 port map( A1 => n1204, A2 => n291, ZN => CU_Ixcw2_6_port);
   U2753 : NOR2_X1 port map( A1 => n1199, A2 => n291, ZN => CU_Ixcw2_1_port);
   U2754 : NOR2_X1 port map( A1 => n1200, A2 => n291, ZN => CU_Ixcw2_2_port);
   U2755 : NOR2_X1 port map( A1 => n1201, A2 => n291, ZN => CU_Ixcw2_3_port);
   U2756 : NOR2_X1 port map( A1 => n1202, A2 => n291, ZN => CU_Ixcw2_4_port);
   U2757 : NOR2_X1 port map( A1 => n1203, A2 => n291, ZN => CU_Ixcw2_5_port);
   U2758 : OR3_X1 port map( A1 => n1411, A2 => n1410, A3 => n144, ZN => n132);
   U2759 : OR3_X1 port map( A1 => n1405, A2 => n1404, A3 => n1972, ZN => n172);
   U2760 : OR3_X1 port map( A1 => n1401, A2 => n1400, A3 => n1973, ZN => n198);
   U2761 : OR3_X1 port map( A1 => n1409, A2 => n1408, A3 => n1971, ZN => n144);
   U2762 : INV_X1 port map( A => IRAM_DOUT(1), ZN => n1799);
   U2763 : INV_X1 port map( A => IRAM_DOUT(0), ZN => n1800);
   U2764 : NOR3_X1 port map( A1 => n1336, A2 => n1335, A3 => n1663, ZN => n334)
                           ;
   U2765 : XNOR2_X1 port map( A => n1361, B => n1386, ZN => n839);
   U2766 : XNOR2_X1 port map( A => n1357, B => n1386, ZN => n855);
   U2767 : XNOR2_X1 port map( A => n1356, B => n1386, ZN => n854);
   U2768 : XNOR2_X1 port map( A => n1360, B => n1386, ZN => n838);
   U2769 : XNOR2_X1 port map( A => n1355, B => n1657, ZN => n852);
   U2770 : XNOR2_X1 port map( A => n1359, B => n1657, ZN => n836);
   U2771 : NOR3_X1 port map( A1 => n1756, A2 => IRAM_DOUT(14), A3 => 
                           IRAM_DOUT(12), ZN => n38);
   U2772 : AOI21_X1 port map( B1 => n1362, B2 => n1363, A => n1386, ZN => n824)
                           ;
   U2773 : AOI21_X1 port map( B1 => n1358, B2 => n1359, A => n1386, ZN => n843)
                           ;
   U2774 : AOI21_X1 port map( B1 => n1354, B2 => n1355, A => n1386, ZN => n860)
                           ;
   U2775 : XNOR2_X1 port map( A => n1358, B => n1658, ZN => n152);
   U2776 : OAI22_X1 port map( A1 => n1276, A2 => n1745, B1 => n1335, B2 => 
                           n1743, ZN => n1286);
   U2777 : XNOR2_X1 port map( A => n1354, B => n1658, ZN => n180);
   U2778 : OAI22_X1 port map( A1 => n1275, A2 => n1745, B1 => n1336, B2 => 
                           n1743, ZN => n1285);
   U2779 : OAI22_X1 port map( A1 => n1298, A2 => n1923, B1 => n1133, B2 => n26,
                           ZN => CU_IxN51);
   U2780 : OAI22_X1 port map( A1 => n1298, A2 => n1923, B1 => n1133, B2 => 
                           n1134, ZN => CU_IxN52);
   U2781 : OAI21_X1 port map( B1 => n1359, B2 => n1358, A => n1386, ZN => n845)
                           ;
   U2782 : OAI21_X1 port map( B1 => n1355, B2 => n1354, A => n1386, ZN => n862)
                           ;
   U2783 : OAI21_X1 port map( B1 => n1363, B2 => n1362, A => n1386, ZN => n826)
                           ;
   U2784 : OAI22_X1 port map( A1 => n1274, A2 => n1745, B1 => n1664, B2 => 
                           n1743, ZN => n1284);
   U2785 : NOR2_X1 port map( A1 => n1197, A2 => n298, ZN => n1133);
   U2786 : XNOR2_X1 port map( A => n1785, B => IRAM_DOUT(13), ZN => n29);
   U2787 : OR2_X1 port map( A1 => n1672, A2 => n1336, ZN => n1636);
   U2788 : NAND2_X1 port map( A1 => n1344, A2 => n1624, ZN => n950);
   U2789 : NOR3_X1 port map( A1 => n1756, A2 => IRAM_DOUT(5), A3 => 
                           IRAM_DOUT(2), ZN => n43);
   U2790 : NAND2_X1 port map( A1 => n950, A2 => n951, ZN => n946);
   U2791 : AND2_X1 port map( A1 => n1382, A2 => n1342, ZN => n801);
   U2792 : INV_X1 port map( A => IRAM_DOUT(14), ZN => n1785);
   U2793 : INV_X1 port map( A => n35, ZN => n1755);
   U2794 : OAI22_X1 port map( A1 => n26, A2 => n1745, B1 => n1743, B2 => n1275,
                           ZN => n35);
   U2795 : INV_X1 port map( A => IRAM_DOUT(12), ZN => n1787);
   U2796 : AOI22_X1 port map( A1 => n37, A2 => n38, B1 => n1745, B2 => n1623, 
                           ZN => n36);
   U2797 : NOR2_X1 port map( A1 => n1796, A2 => n1786, ZN => n37);
   U2798 : INV_X1 port map( A => n25, ZN => n1754);
   U2799 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n1787, ZN 
                           => n22);
   U2800 : OAI22_X1 port map( A1 => n26, A2 => n1745, B1 => n1743, B2 => n1274,
                           ZN => n25);
   U2801 : INV_X1 port map( A => IRAM_DOUT(13), ZN => n1786);
   U2802 : OR2_X1 port map( A1 => n32, A2 => IRAM_DOUT(13), ZN => n23);
   U2803 : INV_X1 port map( A => n1728, ZN => n1721);
   U2804 : INV_X1 port map( A => n1734, ZN => n1733);
   U2805 : INV_X1 port map( A => n1747, ZN => n1744);
   U2806 : INV_X1 port map( A => Rst, ZN => n1745);
   U2807 : INV_X1 port map( A => Rst, ZN => n1746);
   U2808 : INV_X1 port map( A => Rst, ZN => n1747);
   U2809 : NOR2_X1 port map( A1 => n1751, A2 => n1752, ZN => n1750);
   U2810 : OAI22_X1 port map( A1 => CU_IxN25, A2 => n1753, B1 => CU_IxN24, B2 
                           => n1750, ZN => CU_Ixcw_LUT_0_port);
   U2811 : AOI21_X1 port map( B1 => CU_IxN23, B2 => n1751, A => n1753, ZN => 
                           n1748);
   U2812 : NOR2_X1 port map( A1 => n1750, A2 => n1748, ZN => CU_Ixcw_LUT_1_port
                           );
   U2813 : NOR3_X1 port map( A1 => n1753, A2 => CU_IxN25, A3 => CU_IxN23, ZN =>
                           CU_Ixcw_LUT_2_port);
   U2814 : NOR3_X1 port map( A1 => n1753, A2 => CU_IxN23, A3 => n1751, ZN => 
                           CU_Ixcw_LUT_4_port);
   U2815 : OAI21_X1 port map( B1 => CU_IxN24, B2 => n1752, A => CU_IxN25, ZN =>
                           CU_Ixcw_LUT_5_port);
   U2816 : AOI21_X1 port map( B1 => CU_IxN24, B2 => CU_IxN23, A => n1751, ZN =>
                           CU_Ixcw_LUT_7_port);
   U2817 : OAI22_X1 port map( A1 => CU_IxN24, A2 => n1751, B1 => n1750, B2 => 
                           n1753, ZN => CU_Ixcw_LUT_8_port);
   U2818 : NOR2_X1 port map( A1 => CU_IxN24, A2 => CU_IxN25, ZN => 
                           CU_Ixcw_LUT_10_port);
   U2819 : NAND2_X1 port map( A1 => CU_Ixcw_LUT_10_port, A2 => CU_IxN23, ZN => 
                           n1749);
   U2820 : OAI21_X1 port map( B1 => n1751, B2 => n1753, A => n1749, ZN => 
                           CU_Ixcw_LUT_15_port);
   U2821 : NAND2_X1 port map( A1 => CU_IxN24, A2 => n1750, ZN => 
                           CU_Ixcw_LUT_16_port);
   U2822 : AND2_X1 port map( A1 => n1753, A2 => n1750, ZN => CU_Ixcw_LUT_9_port
                           );
   U2823 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_0_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, S => n1741, Z =>
                           n1978);
   U2824 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_2_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_3_port, S => n1742, Z =>
                           n2074);
   U2825 : MUX2_X1 port map( A => n1978, B => n2074, S => n1739, Z => n1979);
   U2826 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_4_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, S => n1742, Z =>
                           n2073);
   U2827 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_6_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, S => n1742, Z =>
                           n2076);
   U2828 : MUX2_X1 port map( A => n2073, B => n2076, S => n1740, Z => n2096);
   U2829 : MUX2_X1 port map( A => n1979, B => n2096, S => n1737, Z => n1980);
   U2830 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_8_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, S => n1742, Z =>
                           n2075);
   U2831 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_10_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, S => n1742, Z 
                           => n1984);
   U2832 : MUX2_X1 port map( A => n2075, B => n1984, S => n1740, Z => n2095);
   U2833 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_12_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, S => n1742, Z 
                           => n1983);
   U2834 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_14_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_15_port, S => n1742, Z 
                           => n1986);
   U2835 : MUX2_X1 port map( A => n1983, B => n1986, S => n1740, Z => n1999);
   U2836 : MUX2_X1 port map( A => n2095, B => n1999, S => n1738, Z => n2124);
   U2837 : MUX2_X1 port map( A => n1980, B => n2124, S => n1735, Z => n1981);
   U2838 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_16_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, S => n1742, Z 
                           => n1985);
   U2839 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_18_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_19_port, S => n1742, Z 
                           => n1988);
   U2840 : MUX2_X1 port map( A => n1985, B => n1988, S => n1740, Z => n1998);
   U2841 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_20_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, S => n1742, Z 
                           => n1987);
   U2842 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_22_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_23_port, S => n1742, Z 
                           => n1990);
   U2843 : MUX2_X1 port map( A => n1987, B => n1990, S => n1740, Z => n2001);
   U2844 : MUX2_X1 port map( A => n1998, B => n2001, S => n1738, Z => n2123);
   U2845 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_24_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, S => n1741, Z 
                           => n1989);
   U2846 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_26_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_27_port, S => n1741, Z 
                           => n1992);
   U2847 : MUX2_X1 port map( A => n1989, B => n1992, S => n1740, Z => n2000);
   U2848 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_28_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, S => n1741, Z 
                           => n1991);
   U2849 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_30_port, B => 
                           n1638, S => n1741, Z => n1993);
   U2850 : MUX2_X1 port map( A => n1991, B => n1993, S => n1740, Z => n2002);
   U2851 : MUX2_X1 port map( A => n2000, B => n2002, S => n1738, Z => n2061);
   U2852 : MUX2_X1 port map( A => n2123, B => n2061, S => n1736, Z => n2029);
   U2853 : MUX2_X1 port map( A => n1981, B => n2029, S => n1733, Z => n1982);
   U2854 : MUX2_X1 port map( A => n1982, B => n1639, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN191);
   U2855 : MUX2_X1 port map( A => n1984, B => n1983, S => n1740, Z => n2109);
   U2856 : MUX2_X1 port map( A => n1986, B => n1985, S => n1740, Z => n2017);
   U2857 : MUX2_X1 port map( A => n2109, B => n2017, S => n1738, Z => n2078);
   U2858 : MUX2_X1 port map( A => n1988, B => n1987, S => n1740, Z => n2016);
   U2859 : MUX2_X1 port map( A => n1990, B => n1989, S => n1740, Z => n2019);
   U2860 : MUX2_X1 port map( A => n2016, B => n2019, S => n1738, Z => n2037);
   U2861 : MUX2_X1 port map( A => n2078, B => n2037, S => n1736, Z => n1994);
   U2862 : MUX2_X1 port map( A => n1992, B => n1991, S => n1739, Z => n2018);
   U2863 : MUX2_X1 port map( A => n1993, B => n1639, S => n1739, Z => n2020);
   U2864 : MUX2_X1 port map( A => n2018, B => n2020, S => n1738, Z => n2036);
   U2865 : MUX2_X1 port map( A => n2036, B => n1639, S => n1736, Z => n2065);
   U2866 : MUX2_X1 port map( A => n1994, B => n2065, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n1995);
   U2867 : MUX2_X1 port map( A => n1995, B => n1639, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN201);
   U2868 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_11_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, S => n1741, Z 
                           => n2044);
   U2869 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_13_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_14_port, S => n1741, Z 
                           => n2006);
   U2870 : MUX2_X1 port map( A => n2044, B => n2006, S => n1739, Z => n2116);
   U2871 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_15_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_16_port, S => n1741, Z 
                           => n2005);
   U2872 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_17_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, S => n1741, Z 
                           => n2008);
   U2873 : MUX2_X1 port map( A => n2005, B => n2008, S => n1739, Z => n2024);
   U2874 : MUX2_X1 port map( A => n2116, B => n2024, S => n1738, Z => n2090);
   U2875 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_19_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, S => n1741, Z 
                           => n2007);
   U2876 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_21_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_22_port, S => n1741, Z 
                           => n2010);
   U2877 : MUX2_X1 port map( A => n2007, B => n2010, S => n1739, Z => n2023);
   U2878 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_23_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, S => n1741, Z 
                           => n2009);
   U2879 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_25_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_26_port, S => n1741, Z 
                           => n2012);
   U2880 : MUX2_X1 port map( A => n2009, B => n2012, S => n1739, Z => n2026);
   U2881 : MUX2_X1 port map( A => n2023, B => n2026, S => n1738, Z => n2040);
   U2882 : MUX2_X1 port map( A => n2090, B => n2040, S => n1736, Z => n1996);
   U2883 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_27_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, S => n1741, Z 
                           => n2011);
   U2884 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_29_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, S => n1741, Z 
                           => n2013);
   U2885 : MUX2_X1 port map( A => n2011, B => n2013, S => n1739, Z => n2025);
   U2886 : MUX2_X1 port map( A => n2025, B => n1639, S => n1738, Z => n2039);
   U2887 : MUX2_X1 port map( A => n2039, B => n1639, S => n1736, Z => n2067);
   U2888 : MUX2_X1 port map( A => n1996, B => n2067, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n1997);
   U2889 : MUX2_X1 port map( A => n1997, B => n1639, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN202);
   U2890 : MUX2_X1 port map( A => n1999, B => n1998, S => n1738, Z => n2097);
   U2891 : MUX2_X1 port map( A => n2001, B => n2000, S => n1738, Z => n2051);
   U2892 : MUX2_X1 port map( A => n2097, B => n2051, S => n1736, Z => n2003);
   U2893 : MUX2_X1 port map( A => n2002, B => n1639, S => n1738, Z => n2050);
   U2894 : MUX2_X1 port map( A => n2050, B => n1639, S => n1736, Z => n2069);
   U2895 : MUX2_X1 port map( A => n2003, B => n2069, S => n1733, Z => n2004);
   U2896 : MUX2_X1 port map( A => n2004, B => n1639, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN203);
   U2897 : MUX2_X1 port map( A => n2006, B => n2005, S => n1739, Z => n2045);
   U2898 : MUX2_X1 port map( A => n2008, B => n2007, S => n1739, Z => n2032);
   U2899 : MUX2_X1 port map( A => n2045, B => n2032, S => n1737, Z => n2104);
   U2900 : MUX2_X1 port map( A => n2010, B => n2009, S => n1739, Z => n2031);
   U2901 : MUX2_X1 port map( A => n2012, B => n2011, S => n1739, Z => n2034);
   U2902 : MUX2_X1 port map( A => n2031, B => n2034, S => n1737, Z => n2054);
   U2903 : MUX2_X1 port map( A => n2104, B => n2054, S => n1736, Z => n2014);
   U2904 : MUX2_X1 port map( A => n2013, B => n1639, S => n1739, Z => n2033);
   U2905 : MUX2_X1 port map( A => n2033, B => n1638, S => n1737, Z => n2053);
   U2906 : MUX2_X1 port map( A => n2053, B => n1638, S => n1736, Z => n2071);
   U2907 : MUX2_X1 port map( A => n2014, B => n2071, S => n1733, Z => n2015);
   U2908 : MUX2_X1 port map( A => n2015, B => n1638, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN204);
   U2909 : MUX2_X1 port map( A => n2017, B => n2016, S => n1737, Z => n2111);
   U2910 : MUX2_X1 port map( A => n2019, B => n2018, S => n1737, Z => n2057);
   U2911 : MUX2_X1 port map( A => n2111, B => n2057, S => n1736, Z => n2021);
   U2912 : MUX2_X1 port map( A => n2020, B => n1638, S => n1737, Z => n2056);
   U2913 : MUX2_X1 port map( A => n2056, B => n1638, S => n1736, Z => n2083);
   U2914 : MUX2_X1 port map( A => n2021, B => n2083, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2022);
   U2915 : MUX2_X1 port map( A => n2022, B => n1638, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN205);
   U2916 : MUX2_X1 port map( A => n2024, B => n2023, S => n1737, Z => n2118);
   U2917 : MUX2_X1 port map( A => n2026, B => n2025, S => n1737, Z => n2059);
   U2918 : MUX2_X1 port map( A => n2118, B => n2059, S => n1736, Z => n2027);
   U2919 : MUX2_X1 port map( A => n2027, B => n1638, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2028);
   U2920 : MUX2_X1 port map( A => n2028, B => n1638, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN206);
   U2921 : MUX2_X1 port map( A => n2029, B => n1638, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2030);
   U2922 : MUX2_X1 port map( A => n2030, B => n1638, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN207);
   U2923 : MUX2_X1 port map( A => n2032, B => n2031, S => n1737, Z => n2128);
   U2924 : MUX2_X1 port map( A => n2034, B => n2033, S => n1737, Z => n2063);
   U2925 : MUX2_X1 port map( A => n2128, B => n2063, S => n1735, Z => n2047);
   U2926 : MUX2_X1 port map( A => n2047, B => n1638, S => n1733, Z => n2035);
   U2927 : MUX2_X1 port map( A => n2035, B => n1637, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN208);
   U2928 : MUX2_X1 port map( A => n2037, B => n2036, S => n1735, Z => n2080);
   U2929 : MUX2_X1 port map( A => n2080, B => n1637, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2038);
   U2930 : MUX2_X1 port map( A => n2038, B => n1637, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN209);
   U2931 : MUX2_X1 port map( A => n2040, B => n2039, S => n1735, Z => n2092);
   U2932 : MUX2_X1 port map( A => n2092, B => n1637, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2041);
   U2933 : MUX2_X1 port map( A => n2041, B => n1637, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN210);
   U2934 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_1_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_2_port, S => n1741, Z =>
                           n2042);
   U2935 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_3_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, S => n1741, Z =>
                           n2086);
   U2936 : MUX2_X1 port map( A => n2042, B => n2086, S => n1739, Z => n2043);
   U2937 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_5_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_6_port, S => n1741, Z =>
                           n2085);
   U2938 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_7_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, S => n1741, Z =>
                           n2088);
   U2939 : MUX2_X1 port map( A => n2085, B => n2088, S => n1739, Z => n2103);
   U2940 : MUX2_X1 port map( A => n2043, B => n2103, S => n1737, Z => n2046);
   U2941 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_9_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, S => n1741, Z 
                           => n2087);
   U2942 : MUX2_X1 port map( A => n2087, B => n2044, S => n1739, Z => n2102);
   U2943 : MUX2_X1 port map( A => n2102, B => n2045, S => n1737, Z => n2129);
   U2944 : MUX2_X1 port map( A => n2046, B => n2129, S => n1735, Z => n2048);
   U2945 : MUX2_X1 port map( A => n2048, B => n2047, S => 
                           DATAPATH_IxThird_stxALU_IN2_4_port, Z => n2049);
   U2946 : MUX2_X1 port map( A => n2049, B => n1637, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN192);
   U2947 : MUX2_X1 port map( A => n2051, B => n2050, S => n1735, Z => n2099);
   U2948 : MUX2_X1 port map( A => n2099, B => n1637, S => n1733, Z => n2052);
   U2949 : MUX2_X1 port map( A => n2052, B => n1637, S => n1730, Z => 
                           DATAPATH_IxThird_stxALU1xN211);
   U2950 : MUX2_X1 port map( A => n2054, B => n2053, S => n1735, Z => n2106);
   U2951 : MUX2_X1 port map( A => n2106, B => n1637, S => n1733, Z => n2055);
   U2952 : MUX2_X1 port map( A => n2055, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN212);
   U2953 : MUX2_X1 port map( A => n2057, B => n2056, S => n1735, Z => n2113);
   U2954 : MUX2_X1 port map( A => n2113, B => n1637, S => n1733, Z => n2058);
   U2955 : MUX2_X1 port map( A => n2058, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN213);
   U2956 : MUX2_X1 port map( A => n2059, B => n1637, S => n1735, Z => n2120);
   U2957 : MUX2_X1 port map( A => n2120, B => n1638, S => n1733, Z => n2060);
   U2958 : MUX2_X1 port map( A => n2060, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN214);
   U2959 : MUX2_X1 port map( A => n2061, B => n1637, S => n1735, Z => n2125);
   U2960 : MUX2_X1 port map( A => n2125, B => n1637, S => n1733, Z => n2062);
   U2961 : MUX2_X1 port map( A => n2062, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN215);
   U2962 : MUX2_X1 port map( A => n2063, B => n1637, S => n1735, Z => n2130);
   U2963 : MUX2_X1 port map( A => n2130, B => n1638, S => n1733, Z => n2064);
   U2964 : MUX2_X1 port map( A => n2064, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN216);
   U2965 : MUX2_X1 port map( A => n2065, B => n1637, S => n1733, Z => n2066);
   U2966 : MUX2_X1 port map( A => n2066, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN217);
   U2967 : MUX2_X1 port map( A => n2067, B => n1637, S => n1733, Z => n2068);
   U2968 : MUX2_X1 port map( A => n2068, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN218);
   U2969 : MUX2_X1 port map( A => n2069, B => n1637, S => n1733, Z => n2070);
   U2970 : MUX2_X1 port map( A => n2070, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN219);
   U2971 : MUX2_X1 port map( A => n2071, B => n1638, S => n1733, Z => n2072);
   U2972 : MUX2_X1 port map( A => n2072, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN220);
   U2973 : MUX2_X1 port map( A => n2074, B => n2073, S => n1739, Z => n2077);
   U2974 : MUX2_X1 port map( A => n2076, B => n2075, S => n1739, Z => n2110);
   U2975 : MUX2_X1 port map( A => n2077, B => n2110, S => n1737, Z => n2079);
   U2976 : MUX2_X1 port map( A => n2079, B => n2078, S => n1735, Z => n2081);
   U2977 : MUX2_X1 port map( A => n2081, B => n2080, S => n1733, Z => n2082);
   U2978 : MUX2_X1 port map( A => n2082, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN193);
   U2979 : MUX2_X1 port map( A => n2083, B => n1638, S => n1733, Z => n2084);
   U2980 : MUX2_X1 port map( A => n2084, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN221);
   U2981 : MUX2_X1 port map( A => n2086, B => n2085, S => n1739, Z => n2089);
   U2982 : MUX2_X1 port map( A => n2088, B => n2087, S => n1739, Z => n2117);
   U2983 : MUX2_X1 port map( A => n2089, B => n2117, S => n1737, Z => n2091);
   U2984 : MUX2_X1 port map( A => n2091, B => n2090, S => n1735, Z => n2093);
   U2985 : MUX2_X1 port map( A => n2093, B => n2092, S => n1733, Z => n2094);
   U2986 : MUX2_X1 port map( A => n2094, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN194);
   U2987 : MUX2_X1 port map( A => n2096, B => n2095, S => n1737, Z => n2098);
   U2988 : MUX2_X1 port map( A => n2098, B => n2097, S => n1735, Z => n2100);
   U2989 : MUX2_X1 port map( A => n2100, B => n2099, S => n1733, Z => n2101);
   U2990 : MUX2_X1 port map( A => n2101, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN195);
   U2991 : MUX2_X1 port map( A => n2103, B => n2102, S => n1737, Z => n2105);
   U2992 : MUX2_X1 port map( A => n2105, B => n2104, S => n1735, Z => n2107);
   U2993 : MUX2_X1 port map( A => n2107, B => n2106, S => n1733, Z => n2108);
   U2994 : MUX2_X1 port map( A => n2108, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN196);
   U2995 : MUX2_X1 port map( A => n2110, B => n2109, S => n1737, Z => n2112);
   U2996 : MUX2_X1 port map( A => n2112, B => n2111, S => n1735, Z => n2114);
   U2997 : MUX2_X1 port map( A => n2114, B => n2113, S => n1733, Z => n2115);
   U2998 : MUX2_X1 port map( A => n2115, B => n1638, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN197);
   U2999 : MUX2_X1 port map( A => n2117, B => n2116, S => n1737, Z => n2119);
   U3000 : MUX2_X1 port map( A => n2119, B => n2118, S => n1735, Z => n2121);
   U3001 : MUX2_X1 port map( A => n2121, B => n2120, S => n1733, Z => n2122);
   U3002 : MUX2_X1 port map( A => n2122, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN198);
   U3003 : MUX2_X1 port map( A => n2124, B => n2123, S => n1735, Z => n2126);
   U3004 : MUX2_X1 port map( A => n2126, B => n2125, S => n1733, Z => n2127);
   U3005 : MUX2_X1 port map( A => n2127, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN199);
   U3006 : MUX2_X1 port map( A => n2129, B => n2128, S => n1735, Z => n2131);
   U3007 : MUX2_X1 port map( A => n2131, B => n2130, S => n1733, Z => n2132);
   U3008 : MUX2_X1 port map( A => n2132, B => n1637, S => n1731, Z => 
                           DATAPATH_IxThird_stxALU1xN200);

end SYN_RV32I_rtl;
