
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RV32I is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RV32I;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RV32I.all;

entity RV32I is

   port( Clk, Rst : in std_logic;  IRAM_DOUT, RF_RD1_DATA, RF_RD2_DATA, 
         DRAM_DOUT : in std_logic_vector (31 downto 0);  IRAM_ADD : out 
         std_logic_vector (31 downto 0);  RF_RD1_EN, RF_RD2_EN, RF_WR_EN : out 
         std_logic;  RF_RD1_ADD, RF_RD2_ADD, RF_WR_ADD : out std_logic_vector 
         (4 downto 0);  RF_WR_DATA : out std_logic_vector (31 downto 0);  
         DRAM_WE, DRAM_RE : out std_logic;  DRAM_ADD, DRAM_DIN : out 
         std_logic_vector (31 downto 0));

end RV32I;

architecture SYN_RV32I_rtl of RV32I is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, RF_RD1_ADD_4_port, 
      RF_RD1_ADD_3_port, RF_RD1_ADD_2_port, RF_RD1_ADD_1_port, 
      RF_RD1_ADD_0_port, RF_RD2_ADD_4_port, RF_RD2_ADD_3_port, 
      RF_RD2_ADD_2_port, RF_RD2_ADD_1_port, RF_RD2_ADD_0_port, n2365, 
      DRAM_ADD_31_port, DRAM_ADD_30_port, DRAM_ADD_29_port, DRAM_ADD_28_port, 
      DRAM_ADD_27_port, DRAM_ADD_26_port, DRAM_ADD_25_port, DRAM_ADD_24_port, 
      DRAM_ADD_23_port, DRAM_ADD_22_port, DRAM_ADD_21_port, DRAM_ADD_20_port, 
      DRAM_ADD_19_port, DRAM_ADD_18_port, DRAM_ADD_17_port, DRAM_ADD_16_port, 
      DRAM_ADD_15_port, DRAM_ADD_14_port, DRAM_ADD_13_port, DRAM_ADD_12_port, 
      DRAM_ADD_11_port, DRAM_ADD_10_port, DRAM_ADD_9_port, DRAM_ADD_8_port, 
      DRAM_ADD_7_port, DRAM_ADD_6_port, DRAM_ADD_5_port, DRAM_ADD_4_port, 
      DRAM_ADD_3_port, DRAM_ADD_2_port, DRAM_ADD_1_port, DRAM_ADD_0_port, 
      PC_SEL_i, IMM_SEL_i, RF_WE_MEM_i, WB_MUX_SEL_MEM_i, BRANCH_EN_i, CU_IxN52
      , CU_IxN51, CU_Ixcw2_i_10_port, CU_Ixcw2_i_11_port, CU_Ixcw2_i_12_port, 
      CU_Ixcw3_0_port, CU_Ixcw3_1_port, CU_Ixcw3_2_port, CU_Ixcw3_3_port, 
      CU_Ixcw2_0_port, CU_Ixcw2_1_port, CU_Ixcw2_2_port, CU_Ixcw2_3_port, 
      CU_Ixcw2_4_port, CU_Ixcw2_5_port, CU_Ixcw2_6_port, CU_Ixcw1_0_port, 
      CU_Ixcw1_1_port, CU_Ixcw1_2_port, CU_Ixcw1_4_port, CU_Ixcw1_5_port, 
      CU_Ixcw1_6_port, CU_Ixcw1_7_port, CU_Ixcw1_8_port, CU_Ixcw1_9_port, 
      CU_Ixcw1_10_port, CU_Ixcw1_14_port, CU_Ixcw_LUT_0_port, 
      CU_Ixcw_LUT_1_port, CU_Ixcw_LUT_2_port, CU_Ixcw_LUT_4_port, 
      CU_Ixcw_LUT_5_port, CU_Ixcw_LUT_6_port, CU_Ixcw_LUT_7_port, 
      CU_Ixcw_LUT_8_port, CU_Ixcw_LUT_9_port, CU_Ixcw_LUT_10_port, 
      CU_Ixcw_LUT_15_port, CU_Ixcw_LUT_16_port, CU_IxN25, CU_IxN24, CU_IxN23, 
      DATAPATH_IxALUOUT_Data1_0_port, DATAPATH_IxALUOUT_Data1_1_port, 
      DATAPATH_IxALUOUT_Data1_2_port, DATAPATH_IxALUOUT_Data1_3_port, 
      DATAPATH_IxALUOUT_Data1_4_port, DATAPATH_IxALUOUT_Data1_5_port, 
      DATAPATH_IxALUOUT_Data1_6_port, DATAPATH_IxALUOUT_Data1_7_port, 
      DATAPATH_IxALUOUT_Data1_8_port, DATAPATH_IxALUOUT_Data1_9_port, 
      DATAPATH_IxALUOUT_Data1_10_port, DATAPATH_IxALUOUT_Data1_11_port, 
      DATAPATH_IxALUOUT_Data1_12_port, DATAPATH_IxALUOUT_Data1_13_port, 
      DATAPATH_IxALUOUT_Data1_14_port, DATAPATH_IxALUOUT_Data1_15_port, 
      DATAPATH_IxALUOUT_Data1_16_port, DATAPATH_IxALUOUT_Data1_17_port, 
      DATAPATH_IxALUOUT_Data1_18_port, DATAPATH_IxALUOUT_Data1_19_port, 
      DATAPATH_IxALUOUT_Data1_20_port, DATAPATH_IxALUOUT_Data1_21_port, 
      DATAPATH_IxALUOUT_Data1_22_port, DATAPATH_IxALUOUT_Data1_23_port, 
      DATAPATH_IxALUOUT_Data1_24_port, DATAPATH_IxALUOUT_Data1_25_port, 
      DATAPATH_IxALUOUT_Data1_26_port, DATAPATH_IxALUOUT_Data1_27_port, 
      DATAPATH_IxALUOUT_Data1_28_port, DATAPATH_IxALUOUT_Data1_29_port, 
      DATAPATH_IxALUOUT_Data1_30_port, DATAPATH_IxALUOUT_Data1_31_port, 
      DATAPATH_IxLMD_DATA_0_port, DATAPATH_IxLMD_DATA_1_port, 
      DATAPATH_IxLMD_DATA_2_port, DATAPATH_IxLMD_DATA_3_port, 
      DATAPATH_IxLMD_DATA_4_port, DATAPATH_IxLMD_DATA_5_port, 
      DATAPATH_IxLMD_DATA_6_port, DATAPATH_IxLMD_DATA_7_port, 
      DATAPATH_IxLMD_DATA_8_port, DATAPATH_IxLMD_DATA_9_port, 
      DATAPATH_IxLMD_DATA_10_port, DATAPATH_IxLMD_DATA_11_port, 
      DATAPATH_IxLMD_DATA_12_port, DATAPATH_IxLMD_DATA_13_port, 
      DATAPATH_IxLMD_DATA_14_port, DATAPATH_IxLMD_DATA_15_port, 
      DATAPATH_IxLMD_DATA_16_port, DATAPATH_IxLMD_DATA_17_port, 
      DATAPATH_IxLMD_DATA_18_port, DATAPATH_IxLMD_DATA_19_port, 
      DATAPATH_IxLMD_DATA_20_port, DATAPATH_IxLMD_DATA_21_port, 
      DATAPATH_IxLMD_DATA_22_port, DATAPATH_IxLMD_DATA_23_port, 
      DATAPATH_IxLMD_DATA_24_port, DATAPATH_IxLMD_DATA_25_port, 
      DATAPATH_IxLMD_DATA_26_port, DATAPATH_IxLMD_DATA_27_port, 
      DATAPATH_IxLMD_DATA_28_port, DATAPATH_IxLMD_DATA_29_port, 
      DATAPATH_IxLMD_DATA_30_port, DATAPATH_IxLMD_DATA_31_port, 
      DATAPATH_IxWR_ADD_MEM_fu_0_port, DATAPATH_IxWR_ADD_MEM_fu_1_port, 
      DATAPATH_IxWR_ADD_MEM_fu_2_port, DATAPATH_IxWR_ADD_MEM_fu_3_port, 
      DATAPATH_IxWR_ADD_MEM_fu_4_port, DATAPATH_IxPC4_0_port, 
      DATAPATH_IxPC4_1_port, DATAPATH_IxINSTR_7_port, DATAPATH_IxINSTR_8_port, 
      DATAPATH_IxINSTR_9_port, DATAPATH_IxINSTR_10_port, 
      DATAPATH_IxINSTR_11_port, DATAPATH_IxSecond_stxWRADD_d1_0_port, 
      DATAPATH_IxSecond_stxWRADD_d1_1_port, 
      DATAPATH_IxSecond_stxWRADD_d1_2_port, 
      DATAPATH_IxSecond_stxWRADD_d1_3_port, 
      DATAPATH_IxSecond_stxWRADD_d1_4_port, 
      DATAPATH_IxSecond_stximm_extended_0_port, 
      DATAPATH_IxSecond_stximm_extended_1_port, 
      DATAPATH_IxSecond_stximm_extended_2_port, 
      DATAPATH_IxSecond_stximm_extended_3_port, 
      DATAPATH_IxSecond_stximm_extended_4_port, 
      DATAPATH_IxSecond_stximm_extended_12_port, 
      DATAPATH_IxSecond_stximm_extended_13_port, 
      DATAPATH_IxSecond_stximm_extended_14_port, 
      DATAPATH_IxSecond_stximm_extended_15_port, 
      DATAPATH_IxSecond_stximm_extended_16_port, 
      DATAPATH_IxSecond_stximm_extended_17_port, 
      DATAPATH_IxSecond_stximm_extended_18_port, 
      DATAPATH_IxSecond_stximm_extended_19_port, 
      DATAPATH_IxSecond_stximm_extended_20_port, 
      DATAPATH_IxSecond_stximm_extended_21_port, 
      DATAPATH_IxSecond_stximm_extended_22_port, 
      DATAPATH_IxSecond_stximm_extended_23_port, 
      DATAPATH_IxSecond_stximm_extended_24_port, 
      DATAPATH_IxSecond_stximm_extended_25_port, 
      DATAPATH_IxSecond_stximm_extended_26_port, 
      DATAPATH_IxSecond_stximm_extended_27_port, 
      DATAPATH_IxSecond_stximm_extended_28_port, 
      DATAPATH_IxSecond_stximm_extended_29_port, 
      DATAPATH_IxSecond_stximm_extended_30_port, 
      DATAPATH_IxSecond_stximm_extended_31_port, 
      DATAPATH_IxSecond_stxBR_target_2_port, 
      DATAPATH_IxSecond_stxBR_target_6_port, 
      DATAPATH_IxSecond_stxBR_target_8_port, 
      DATAPATH_IxSecond_stxBR_target_10_port, 
      DATAPATH_IxSecond_stxBR_target_12_port, 
      DATAPATH_IxSecond_stxBR_target_14_port, 
      DATAPATH_IxSecond_stxBR_target_18_port, 
      DATAPATH_IxSecond_stxjump_target_0_port, 
      DATAPATH_IxSecond_stxjump_target_3_port, 
      DATAPATH_IxSecond_stxjump_target_5_port, 
      DATAPATH_IxSecond_stxjump_target_6_port, 
      DATAPATH_IxSecond_stxjump_target_7_port, 
      DATAPATH_IxSecond_stxjump_target_10_port, 
      DATAPATH_IxSecond_stxjump_target_11_port, 
      DATAPATH_IxSecond_stxjump_target_12_port, 
      DATAPATH_IxSecond_stxjump_target_14_port, 
      DATAPATH_IxSecond_stxjump_target_16_port, 
      DATAPATH_IxSecond_stxjump_target_17_port, 
      DATAPATH_IxSecond_stxjump_target_18_port, 
      DATAPATH_IxSecond_stxjump_target_21_port, 
      DATAPATH_IxSecond_stxjump_target_22_port, 
      DATAPATH_IxSecond_stxjump_target_23_port, 
      DATAPATH_IxSecond_stxjump_target_25_port, 
      DATAPATH_IxSecond_stxjump_target_26_port, 
      DATAPATH_IxSecond_stxjump_target_27_port, 
      DATAPATH_IxSecond_stxjump_target_30_port, 
      DATAPATH_IxSecond_stxjump_target_31_port, 
      DATAPATH_IxThird_stxALU_out_i_0_port, 
      DATAPATH_IxThird_stxALU_out_i_1_port, 
      DATAPATH_IxThird_stxALU_out_i_2_port, 
      DATAPATH_IxThird_stxALU_out_i_3_port, 
      DATAPATH_IxThird_stxALU_out_i_4_port, 
      DATAPATH_IxThird_stxALU_out_i_5_port, 
      DATAPATH_IxThird_stxALU_out_i_6_port, 
      DATAPATH_IxThird_stxALU_out_i_7_port, 
      DATAPATH_IxThird_stxALU_out_i_8_port, 
      DATAPATH_IxThird_stxALU_out_i_9_port, 
      DATAPATH_IxThird_stxALU_out_i_10_port, 
      DATAPATH_IxThird_stxALU_out_i_11_port, 
      DATAPATH_IxThird_stxALU_out_i_12_port, 
      DATAPATH_IxThird_stxALU_out_i_13_port, 
      DATAPATH_IxThird_stxALU_out_i_14_port, 
      DATAPATH_IxThird_stxALU_out_i_15_port, 
      DATAPATH_IxThird_stxALU_out_i_16_port, 
      DATAPATH_IxThird_stxALU_out_i_17_port, 
      DATAPATH_IxThird_stxALU_out_i_18_port, 
      DATAPATH_IxThird_stxALU_out_i_19_port, 
      DATAPATH_IxThird_stxALU_out_i_20_port, 
      DATAPATH_IxThird_stxALU_out_i_21_port, 
      DATAPATH_IxThird_stxALU_out_i_22_port, 
      DATAPATH_IxThird_stxALU_out_i_23_port, 
      DATAPATH_IxThird_stxALU_out_i_24_port, 
      DATAPATH_IxThird_stxALU_out_i_25_port, 
      DATAPATH_IxThird_stxALU_out_i_26_port, 
      DATAPATH_IxThird_stxALU_out_i_27_port, 
      DATAPATH_IxThird_stxALU_out_i_28_port, 
      DATAPATH_IxThird_stxALU_out_i_29_port, 
      DATAPATH_IxThird_stxALU_out_i_30_port, 
      DATAPATH_IxThird_stxALU_out_i_31_port, DATAPATH_IxThird_stxALU_IN2_0_port
      , DATAPATH_IxThird_stxALU_IN2_1_port, DATAPATH_IxThird_stxALU_IN2_2_port,
      DATAPATH_IxThird_stxALU_IN2_3_port, DATAPATH_IxThird_stxALU_IN2_4_port, 
      DATAPATH_IxThird_stxALU_IN2_5_port, DATAPATH_IxThird_stxALU_IN1_0_port, 
      DATAPATH_IxThird_stxALU_IN1_1_port, DATAPATH_IxThird_stxALU_IN1_2_port, 
      DATAPATH_IxThird_stxALU_IN1_3_port, DATAPATH_IxThird_stxALU_IN1_4_port, 
      DATAPATH_IxThird_stxALU_IN1_5_port, DATAPATH_IxThird_stxALU_IN1_6_port, 
      DATAPATH_IxThird_stxALU_IN1_7_port, DATAPATH_IxThird_stxALU_IN1_8_port, 
      DATAPATH_IxThird_stxALU_IN1_9_port, DATAPATH_IxThird_stxALU_IN1_10_port, 
      DATAPATH_IxThird_stxALU_IN1_11_port, DATAPATH_IxThird_stxALU_IN1_12_port,
      DATAPATH_IxThird_stxALU_IN1_13_port, DATAPATH_IxThird_stxALU_IN1_14_port,
      DATAPATH_IxThird_stxALU_IN1_15_port, DATAPATH_IxThird_stxALU_IN1_16_port,
      DATAPATH_IxThird_stxALU_IN1_17_port, DATAPATH_IxThird_stxALU_IN1_18_port,
      DATAPATH_IxThird_stxALU_IN1_19_port, DATAPATH_IxThird_stxALU_IN1_20_port,
      DATAPATH_IxThird_stxALU_IN1_21_port, DATAPATH_IxThird_stxALU_IN1_22_port,
      DATAPATH_IxThird_stxALU_IN1_23_port, DATAPATH_IxThird_stxALU_IN1_24_port,
      DATAPATH_IxThird_stxALU_IN1_25_port, DATAPATH_IxThird_stxALU_IN1_26_port,
      DATAPATH_IxThird_stxALU_IN1_27_port, DATAPATH_IxThird_stxALU_IN1_28_port,
      DATAPATH_IxThird_stxALU_IN1_29_port, DATAPATH_IxThird_stxALU_IN1_30_port,
      DATAPATH_IxThird_stxALU1xN222, DATAPATH_IxThird_stxALU1xN221, 
      DATAPATH_IxThird_stxALU1xN220, DATAPATH_IxThird_stxALU1xN219, 
      DATAPATH_IxThird_stxALU1xN218, DATAPATH_IxThird_stxALU1xN217, 
      DATAPATH_IxThird_stxALU1xN216, DATAPATH_IxThird_stxALU1xN215, 
      DATAPATH_IxThird_stxALU1xN214, DATAPATH_IxThird_stxALU1xN213, 
      DATAPATH_IxThird_stxALU1xN212, DATAPATH_IxThird_stxALU1xN211, 
      DATAPATH_IxThird_stxALU1xN210, DATAPATH_IxThird_stxALU1xN209, 
      DATAPATH_IxThird_stxALU1xN208, DATAPATH_IxThird_stxALU1xN207, 
      DATAPATH_IxThird_stxALU1xN206, DATAPATH_IxThird_stxALU1xN205, 
      DATAPATH_IxThird_stxALU1xN204, DATAPATH_IxThird_stxALU1xN203, 
      DATAPATH_IxThird_stxALU1xN202, DATAPATH_IxThird_stxALU1xN201, 
      DATAPATH_IxThird_stxALU1xN200, DATAPATH_IxThird_stxALU1xN199, 
      DATAPATH_IxThird_stxALU1xN198, DATAPATH_IxThird_stxALU1xN197, 
      DATAPATH_IxThird_stxALU1xN196, DATAPATH_IxThird_stxALU1xN195, 
      DATAPATH_IxThird_stxALU1xN194, DATAPATH_IxThird_stxALU1xN193, 
      DATAPATH_IxThird_stxALU1xN192, DATAPATH_IxThird_stxALU1xN191, n22, n23, 
      n25, n26, n27, n28, n29, n32, n33, n35, n36, n37, n38, n43, n46, n47, n48
      , n49, n54, n91, n92, n96, n97, n99, n101, n103, n105, n106, n108, n109, 
      n110, n111, n112, n113, n115, n118, n119, n120, n122, n124, n129, n130, 
      n132, n134, n135, n137, n139, n141, n143, n144, n145, n146, n148, n150, 
      n152, n154, n156, n158, n159, n160, n161, n162, n164, n165, n167, n168, 
      n169, n171, n172, n174, n175, n177, n179, n180, n181, n182, n183, n185, 
      n187, n188, n189, n190, n191, n192, n194, n196, n197, n198, n200, n201, 
      n203, n205, n206, n207, n209, n211, n212, n213, n214, n216, n217, n218, 
      n219, n221, n222, n223, n224, n226, n228, n229, n231, n232, n233, n234, 
      n236, n237, n238, n239, n241, n242, n243, n244, n246, n248, n250, n251, 
      n253, n254, n255, n256, n258, n260, n261, n262, n265, n266, n267, n268, 
      n269, n270, n271, n273, n275, n278, n279, n280, n282, n283, n284, n285, 
      n286, n289, n291, n292, n294, n296, n298, n299, n326, n328, n330, n331, 
      n333, n334, n335, n336, n337, n338, n340, n344, n345, n346, n347, n348, 
      n349, n351, n352, n353, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n367, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n382, n383, n384, n385, n386, n387, n388, n390, 
      n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n411, n412, n413, n416, n418, n419, n420, n421, 
      n422, n423, n425, n426, n427, n428, n429, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n446, n447, n449, 
      n450, n451, n452, n453, n454, n455, n457, n459, n460, n461, n463, n464, 
      n465, n467, n468, n469, n470, n471, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n483, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n495, n496, n497, n498, n500, n501, n502, n503, n504, n505, n507, 
      n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n532, n534, n535, n536, 
      n537, n538, n539, n540, n541, n543, n544, n545, n546, n548, n549, n550, 
      n551, n552, n553, n555, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n567, n568, n569, n570, n571, n572, n574, n575, n576, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n590, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n605, n607, n608, 
      n609, n610, n611, n613, n615, n616, n617, n618, n619, n620, n622, n623, 
      n624, n625, n626, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n638, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n652, n653, n654, n655, n656, n657, n658, n660, n661, n662, n663, n664, 
      n665, n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n682, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n695, n696, n698, n699, n702, n703, n705, n706, n707, n708, n709, 
      n710, n712, n713, n715, n716, n717, n718, n719, n722, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n737, n738, n739, n740, 
      n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, n753, n754, 
      n755, n757, n758, n759, n760, n762, n765, n766, n767, n768, n769, n770, 
      n771, n773, n774, n775, n776, n778, n779, n780, n781, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n794, n795, n797, n798, n799, 
      n800, n801, n803, n804, n805, n806, n807, n808, n809, n811, n812, n813, 
      n814, n815, n817, n818, n819, n820, n821, n822, n824, n825, n826, n827, 
      n828, n829, n830, n831, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n857, n858, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n876, n877, n878, n879, n882, 
      n884, n885, n886, n887, n889, n890, n894, n896, n897, n898, n899, n900, 
      n901, n903, n904, n905, n906, n907, n909, n910, n911, n912, n913, n914, 
      n915, n916, n917, n918, n919, n920, n921, n922, n924, n925, n927, n929, 
      n930, n931, n932, n933, n934, n936, n938, n939, n940, n941, n942, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n956, n958, 
      n959, n961, n962, n963, n965, n967, n968, n969, n970, n976, n977, n979, 
      n980, n981, n983, n985, n986, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1088, n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1109, n1111, n1113, n1114, n1115, 
      n1116, n1118, n1119, n1120, n1121, n1124, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139, n1140, 
      n1141, n1145, n1146, n1147, n1148, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1241, 
      n1244, n1248, n1257, n1274, n1275, n1276, n1284, n1285, n1286, n1287, 
      n1288, n1289, n1291, n1292, n1296, n1298, n1299, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, RF_WR_DATAx0x, RF_WR_DATAx1x, 
      RF_WR_DATAx2x, RF_WR_DATAx3x, RF_WR_DATAx4x, RF_WR_DATAx5x, RF_WR_DATAx6x
      , RF_WR_DATAx7x, RF_WR_DATAx8x, RF_WR_DATAx9x, RF_WR_DATAx10x, 
      RF_WR_DATAx11x, RF_WR_DATAx12x, RF_WR_DATAx13x, RF_WR_DATAx14x, 
      RF_WR_DATAx15x, RF_WR_DATAx16x, RF_WR_DATAx17x, RF_WR_DATAx18x, 
      RF_WR_DATAx19x, RF_WR_DATAx20x, RF_WR_DATAx21x, RF_WR_DATAx22x, 
      RF_WR_DATAx23x, RF_WR_DATAx24x, RF_WR_DATAx25x, RF_WR_DATAx26x, 
      RF_WR_DATAx27x, RF_WR_DATAx28x, RF_WR_DATAx29x, RF_WR_DATAx30x, 
      RF_WR_DATAx31x, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254 : std_logic;

begin
   IRAM_ADD <= ( IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, DATAPATH_IxPC4_1_port,
      DATAPATH_IxPC4_0_port );
   RF_RD1_ADD <= ( RF_RD1_ADD_4_port, RF_RD1_ADD_3_port, RF_RD1_ADD_2_port, 
      RF_RD1_ADD_1_port, RF_RD1_ADD_0_port );
   RF_RD2_ADD <= ( RF_RD2_ADD_4_port, RF_RD2_ADD_3_port, RF_RD2_ADD_2_port, 
      RF_RD2_ADD_1_port, RF_RD2_ADD_0_port );
   RF_WR_DATA <= ( RF_WR_DATAx31x, RF_WR_DATAx30x, RF_WR_DATAx29x, 
      RF_WR_DATAx28x, RF_WR_DATAx27x, RF_WR_DATAx26x, RF_WR_DATAx25x, 
      RF_WR_DATAx24x, RF_WR_DATAx23x, RF_WR_DATAx22x, RF_WR_DATAx21x, 
      RF_WR_DATAx20x, RF_WR_DATAx19x, RF_WR_DATAx18x, RF_WR_DATAx17x, 
      RF_WR_DATAx16x, RF_WR_DATAx15x, RF_WR_DATAx14x, RF_WR_DATAx13x, 
      RF_WR_DATAx12x, RF_WR_DATAx11x, RF_WR_DATAx10x, RF_WR_DATAx9x, 
      RF_WR_DATAx8x, RF_WR_DATAx7x, RF_WR_DATAx6x, RF_WR_DATAx5x, RF_WR_DATAx4x
      , RF_WR_DATAx3x, RF_WR_DATAx2x, RF_WR_DATAx1x, RF_WR_DATAx0x );
   DRAM_ADD <= ( DRAM_ADD_31_port, DRAM_ADD_30_port, DRAM_ADD_29_port, 
      DRAM_ADD_28_port, DRAM_ADD_27_port, DRAM_ADD_26_port, DRAM_ADD_25_port, 
      DRAM_ADD_24_port, DRAM_ADD_23_port, DRAM_ADD_22_port, DRAM_ADD_21_port, 
      DRAM_ADD_20_port, DRAM_ADD_19_port, DRAM_ADD_18_port, DRAM_ADD_17_port, 
      DRAM_ADD_16_port, DRAM_ADD_15_port, DRAM_ADD_14_port, DRAM_ADD_13_port, 
      DRAM_ADD_12_port, DRAM_ADD_11_port, DRAM_ADD_10_port, DRAM_ADD_9_port, 
      DRAM_ADD_8_port, DRAM_ADD_7_port, DRAM_ADD_6_port, DRAM_ADD_5_port, 
      DRAM_ADD_4_port, DRAM_ADD_3_port, DRAM_ADD_2_port, DRAM_ADD_1_port, 
      DRAM_ADD_0_port );
   
   CU_Ixstate_var_regx1x : DFFR_X1 port map( D => CU_IxN52, CK => Clk, RN => 
                           n1992, Q => n1706, QN => n1197);
   CU_Ixstate_var_regx0x : DFFR_X1 port map( D => CU_IxN51, CK => Clk, RN => 
                           n1991, Q => n1781, QN => n1298);
   CU_IxaluOpcode2_regx0x : DFF_X1 port map( D => n1289, CK => Clk, Q => n1642,
                           QN => n1276);
   CU_IxaluOpcode2_regx1x : DFF_X1 port map( D => n1288, CK => Clk, Q => n_1000
                           , QN => n1275);
   CU_IxaluOpcode2_regx2x : DFF_X1 port map( D => n1287, CK => Clk, Q => n_1001
                           , QN => n1274);
   CU_IxaluOpcode3_regx0x : DFF_X1 port map( D => n1286, CK => Clk, Q => n_1002
                           , QN => n1335);
   CU_IxaluOpcode3_regx1x : DFF_X1 port map( D => n1285, CK => Clk, Q => n1605,
                           QN => n1336);
   CU_IxaluOpcode3_regx2x : DFF_X1 port map( D => n1284, CK => Clk, Q => n1601,
                           QN => n1337);
   DATAPATH_IxThird_stxB_FORWARD_out_regx0x : DFF_X1 port map( D => 
                           RF_RD2_DATA(0), CK => Clk, Q => DRAM_DIN(0), QN => 
                           n_1003);
   DATAPATH_IxThird_stxB_FORWARD_out_regx1x : DFF_X1 port map( D => 
                           RF_RD2_DATA(1), CK => Clk, Q => DRAM_DIN(1), QN => 
                           n_1004);
   DATAPATH_IxThird_stxB_FORWARD_out_regx2x : DFF_X1 port map( D => 
                           RF_RD2_DATA(2), CK => Clk, Q => DRAM_DIN(2), QN => 
                           n_1005);
   DATAPATH_IxThird_stxB_FORWARD_out_regx3x : DFF_X1 port map( D => 
                           RF_RD2_DATA(3), CK => Clk, Q => DRAM_DIN(3), QN => 
                           n_1006);
   DATAPATH_IxThird_stxB_FORWARD_out_regx4x : DFF_X1 port map( D => 
                           RF_RD2_DATA(4), CK => Clk, Q => DRAM_DIN(4), QN => 
                           n_1007);
   DATAPATH_IxThird_stxB_FORWARD_out_regx5x : DFF_X1 port map( D => 
                           RF_RD2_DATA(5), CK => Clk, Q => DRAM_DIN(5), QN => 
                           n_1008);
   DATAPATH_IxThird_stxB_FORWARD_out_regx6x : DFF_X1 port map( D => 
                           RF_RD2_DATA(6), CK => Clk, Q => DRAM_DIN(6), QN => 
                           n_1009);
   DATAPATH_IxThird_stxB_FORWARD_out_regx7x : DFF_X1 port map( D => 
                           RF_RD2_DATA(7), CK => Clk, Q => DRAM_DIN(7), QN => 
                           n_1010);
   DATAPATH_IxThird_stxB_FORWARD_out_regx8x : DFF_X1 port map( D => 
                           RF_RD2_DATA(8), CK => Clk, Q => DRAM_DIN(8), QN => 
                           n_1011);
   DATAPATH_IxThird_stxB_FORWARD_out_regx9x : DFF_X1 port map( D => 
                           RF_RD2_DATA(9), CK => Clk, Q => DRAM_DIN(9), QN => 
                           n_1012);
   DATAPATH_IxThird_stxB_FORWARD_out_regx10x : DFF_X1 port map( D => 
                           RF_RD2_DATA(10), CK => Clk, Q => DRAM_DIN(10), QN =>
                           n_1013);
   DATAPATH_IxThird_stxB_FORWARD_out_regx11x : DFF_X1 port map( D => 
                           RF_RD2_DATA(11), CK => Clk, Q => DRAM_DIN(11), QN =>
                           n_1014);
   DATAPATH_IxThird_stxB_FORWARD_out_regx12x : DFF_X1 port map( D => 
                           RF_RD2_DATA(12), CK => Clk, Q => DRAM_DIN(12), QN =>
                           n_1015);
   DATAPATH_IxThird_stxB_FORWARD_out_regx13x : DFF_X1 port map( D => 
                           RF_RD2_DATA(13), CK => Clk, Q => DRAM_DIN(13), QN =>
                           n_1016);
   DATAPATH_IxThird_stxB_FORWARD_out_regx14x : DFF_X1 port map( D => 
                           RF_RD2_DATA(14), CK => Clk, Q => DRAM_DIN(14), QN =>
                           n_1017);
   DATAPATH_IxThird_stxB_FORWARD_out_regx15x : DFF_X1 port map( D => 
                           RF_RD2_DATA(15), CK => Clk, Q => DRAM_DIN(15), QN =>
                           n_1018);
   DATAPATH_IxThird_stxB_FORWARD_out_regx16x : DFF_X1 port map( D => 
                           RF_RD2_DATA(16), CK => Clk, Q => DRAM_DIN(16), QN =>
                           n_1019);
   DATAPATH_IxThird_stxB_FORWARD_out_regx17x : DFF_X1 port map( D => 
                           RF_RD2_DATA(17), CK => Clk, Q => DRAM_DIN(17), QN =>
                           n_1020);
   DATAPATH_IxThird_stxB_FORWARD_out_regx18x : DFF_X1 port map( D => 
                           RF_RD2_DATA(18), CK => Clk, Q => DRAM_DIN(18), QN =>
                           n_1021);
   DATAPATH_IxThird_stxB_FORWARD_out_regx19x : DFF_X1 port map( D => 
                           RF_RD2_DATA(19), CK => Clk, Q => DRAM_DIN(19), QN =>
                           n_1022);
   DATAPATH_IxThird_stxB_FORWARD_out_regx20x : DFF_X1 port map( D => 
                           RF_RD2_DATA(20), CK => Clk, Q => DRAM_DIN(20), QN =>
                           n_1023);
   DATAPATH_IxThird_stxB_FORWARD_out_regx21x : DFF_X1 port map( D => 
                           RF_RD2_DATA(21), CK => Clk, Q => DRAM_DIN(21), QN =>
                           n_1024);
   DATAPATH_IxThird_stxB_FORWARD_out_regx22x : DFF_X1 port map( D => 
                           RF_RD2_DATA(22), CK => Clk, Q => DRAM_DIN(22), QN =>
                           n_1025);
   DATAPATH_IxThird_stxB_FORWARD_out_regx23x : DFF_X1 port map( D => 
                           RF_RD2_DATA(23), CK => Clk, Q => DRAM_DIN(23), QN =>
                           n_1026);
   DATAPATH_IxThird_stxB_FORWARD_out_regx24x : DFF_X1 port map( D => 
                           RF_RD2_DATA(24), CK => Clk, Q => DRAM_DIN(24), QN =>
                           n_1027);
   DATAPATH_IxThird_stxB_FORWARD_out_regx25x : DFF_X1 port map( D => 
                           RF_RD2_DATA(25), CK => Clk, Q => DRAM_DIN(25), QN =>
                           n_1028);
   DATAPATH_IxThird_stxB_FORWARD_out_regx26x : DFF_X1 port map( D => 
                           RF_RD2_DATA(26), CK => Clk, Q => DRAM_DIN(26), QN =>
                           n_1029);
   DATAPATH_IxThird_stxB_FORWARD_out_regx27x : DFF_X1 port map( D => 
                           RF_RD2_DATA(27), CK => Clk, Q => DRAM_DIN(27), QN =>
                           n_1030);
   DATAPATH_IxThird_stxB_FORWARD_out_regx28x : DFF_X1 port map( D => 
                           RF_RD2_DATA(28), CK => Clk, Q => DRAM_DIN(28), QN =>
                           n_1031);
   DATAPATH_IxThird_stxB_FORWARD_out_regx29x : DFF_X1 port map( D => 
                           RF_RD2_DATA(29), CK => Clk, Q => DRAM_DIN(29), QN =>
                           n_1032);
   DATAPATH_IxThird_stxB_FORWARD_out_regx30x : DFF_X1 port map( D => 
                           RF_RD2_DATA(30), CK => Clk, Q => DRAM_DIN(30), QN =>
                           n_1033);
   DATAPATH_IxThird_stxB_FORWARD_out_regx31x : DFF_X1 port map( D => 
                           RF_RD2_DATA(31), CK => Clk, Q => DRAM_DIN(31), QN =>
                           n_1034);
   DATAPATH_IxFourth_stxLMD_out_regx0x : DFF_X1 port map( D => DRAM_DOUT(0), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_0_port, QN => 
                           n_1035);
   DATAPATH_IxFourth_stxLMD_out_regx1x : DFF_X1 port map( D => DRAM_DOUT(1), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_1_port, QN => 
                           n_1036);
   DATAPATH_IxFourth_stxLMD_out_regx2x : DFF_X1 port map( D => DRAM_DOUT(2), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_2_port, QN => 
                           n_1037);
   DATAPATH_IxFourth_stxLMD_out_regx3x : DFF_X1 port map( D => DRAM_DOUT(3), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_3_port, QN => 
                           n_1038);
   DATAPATH_IxFourth_stxLMD_out_regx4x : DFF_X1 port map( D => DRAM_DOUT(4), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_4_port, QN => 
                           n_1039);
   DATAPATH_IxFourth_stxLMD_out_regx5x : DFF_X1 port map( D => DRAM_DOUT(5), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_5_port, QN => 
                           n_1040);
   DATAPATH_IxFourth_stxLMD_out_regx6x : DFF_X1 port map( D => DRAM_DOUT(6), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_6_port, QN => 
                           n_1041);
   DATAPATH_IxFourth_stxLMD_out_regx7x : DFF_X1 port map( D => DRAM_DOUT(7), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_7_port, QN => 
                           n_1042);
   DATAPATH_IxFourth_stxLMD_out_regx8x : DFF_X1 port map( D => DRAM_DOUT(8), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_8_port, QN => 
                           n_1043);
   DATAPATH_IxFourth_stxLMD_out_regx9x : DFF_X1 port map( D => DRAM_DOUT(9), CK
                           => Clk, Q => DATAPATH_IxLMD_DATA_9_port, QN => 
                           n_1044);
   DATAPATH_IxFourth_stxLMD_out_regx10x : DFF_X1 port map( D => DRAM_DOUT(10), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_10_port, QN => 
                           n_1045);
   DATAPATH_IxFourth_stxLMD_out_regx11x : DFF_X1 port map( D => DRAM_DOUT(11), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_11_port, QN => 
                           n_1046);
   DATAPATH_IxFourth_stxLMD_out_regx12x : DFF_X1 port map( D => DRAM_DOUT(12), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_12_port, QN => 
                           n_1047);
   DATAPATH_IxFourth_stxLMD_out_regx13x : DFF_X1 port map( D => DRAM_DOUT(13), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_13_port, QN => 
                           n_1048);
   DATAPATH_IxFourth_stxLMD_out_regx14x : DFF_X1 port map( D => DRAM_DOUT(14), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_14_port, QN => 
                           n_1049);
   DATAPATH_IxFourth_stxLMD_out_regx15x : DFF_X1 port map( D => DRAM_DOUT(15), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_15_port, QN => 
                           n_1050);
   DATAPATH_IxFourth_stxLMD_out_regx16x : DFF_X1 port map( D => DRAM_DOUT(16), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_16_port, QN => 
                           n_1051);
   DATAPATH_IxFourth_stxLMD_out_regx17x : DFF_X1 port map( D => DRAM_DOUT(17), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_17_port, QN => 
                           n_1052);
   DATAPATH_IxFourth_stxLMD_out_regx18x : DFF_X1 port map( D => DRAM_DOUT(18), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_18_port, QN => 
                           n_1053);
   DATAPATH_IxFourth_stxLMD_out_regx19x : DFF_X1 port map( D => DRAM_DOUT(19), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_19_port, QN => 
                           n_1054);
   DATAPATH_IxFourth_stxLMD_out_regx20x : DFF_X1 port map( D => DRAM_DOUT(20), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_20_port, QN => 
                           n_1055);
   DATAPATH_IxFourth_stxLMD_out_regx21x : DFF_X1 port map( D => DRAM_DOUT(21), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_21_port, QN => 
                           n_1056);
   DATAPATH_IxFourth_stxLMD_out_regx22x : DFF_X1 port map( D => DRAM_DOUT(22), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_22_port, QN => 
                           n_1057);
   DATAPATH_IxFourth_stxLMD_out_regx23x : DFF_X1 port map( D => DRAM_DOUT(23), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_23_port, QN => 
                           n_1058);
   DATAPATH_IxFourth_stxLMD_out_regx24x : DFF_X1 port map( D => DRAM_DOUT(24), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_24_port, QN => 
                           n_1059);
   DATAPATH_IxFourth_stxLMD_out_regx25x : DFF_X1 port map( D => DRAM_DOUT(25), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_25_port, QN => 
                           n_1060);
   DATAPATH_IxFourth_stxLMD_out_regx26x : DFF_X1 port map( D => DRAM_DOUT(26), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_26_port, QN => 
                           n_1061);
   DATAPATH_IxFourth_stxLMD_out_regx27x : DFF_X1 port map( D => DRAM_DOUT(27), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_27_port, QN => 
                           n_1062);
   DATAPATH_IxFourth_stxLMD_out_regx28x : DFF_X1 port map( D => DRAM_DOUT(28), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_28_port, QN => 
                           n_1063);
   DATAPATH_IxFourth_stxLMD_out_regx29x : DFF_X1 port map( D => DRAM_DOUT(29), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_29_port, QN => 
                           n_1064);
   DATAPATH_IxFourth_stxLMD_out_regx30x : DFF_X1 port map( D => DRAM_DOUT(30), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_30_port, QN => 
                           n_1065);
   DATAPATH_IxFourth_stxLMD_out_regx31x : DFF_X1 port map( D => DRAM_DOUT(31), 
                           CK => Clk, Q => DATAPATH_IxLMD_DATA_31_port, QN => 
                           n_1066);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx0x : DFF_X1 port map( D => 
                           DRAM_ADD_0_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_0_port, QN => n_1067);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx10x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_10_port, CK => Clk, Q 
                           => DRAM_ADD_10_port, QN => n1429);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx10x : DFF_X1 port map( D => 
                           DRAM_ADD_10_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_10_port, QN => n_1068);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_16_port, CK => Clk, Q 
                           => DRAM_ADD_16_port, QN => n1435);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx16x : DFF_X1 port map( D => 
                           DRAM_ADD_16_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_16_port, QN => n_1069);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_17_port, CK => Clk, Q 
                           => DRAM_ADD_17_port, QN => n1436);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx17x : DFF_X1 port map( D => 
                           DRAM_ADD_17_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_17_port, QN => n_1070);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_18_port, CK => Clk, Q 
                           => DRAM_ADD_18_port, QN => n1437);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx18x : DFF_X1 port map( D => 
                           DRAM_ADD_18_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_18_port, QN => n_1071);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_25_port, CK => Clk, Q 
                           => DRAM_ADD_25_port, QN => n1444);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx25x : DFF_X1 port map( D => 
                           DRAM_ADD_25_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_25_port, QN => n_1072);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_26_port, CK => Clk, Q 
                           => DRAM_ADD_26_port, QN => n1445);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx26x : DFF_X1 port map( D => 
                           DRAM_ADD_26_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_26_port, QN => n_1073);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_31_port, CK => Clk, Q 
                           => DRAM_ADD_31_port, QN => n1450);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx31x : DFF_X1 port map( D => 
                           DRAM_ADD_31_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_31_port, QN => n_1074);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx31x : DFF_X1 port map( D => n1548, CK 
                           => Clk, Q => n1689, QN => n1386);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx30x : DFF_X1 port map( D => n1549, CK 
                           => Clk, Q => n_1075, QN => n1385);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx29x : DFF_X1 port map( D => n1550, CK 
                           => Clk, Q => n_1076, QN => n1646);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx28x : DFF_X1 port map( D => n1551, CK 
                           => Clk, Q => n_1077, QN => n1384);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx27x : DFF_X1 port map( D => n1552, CK 
                           => Clk, Q => n_1078, QN => n1383);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx26x : DFF_X1 port map( D => n1553, CK 
                           => Clk, Q => n_1079, QN => n1382);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx25x : DFF_X1 port map( D => n1554, CK 
                           => Clk, Q => n_1080, QN => n1381);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx24x : DFF_X1 port map( D => n1555, CK 
                           => Clk, Q => RF_RD2_ADD_4_port, QN => n1380);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx4x : DFF_X1 port map( D => 
                           RF_RD2_ADD_4_port, CK => Clk, Q => n_1081, QN => 
                           n1154);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx23x : DFF_X1 port map( D => n1556, CK 
                           => Clk, Q => RF_RD2_ADD_3_port, QN => n1379);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx22x : DFF_X1 port map( D => n1557, CK 
                           => Clk, Q => RF_RD2_ADD_2_port, QN => n1378);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx2x : DFF_X1 port map( D => 
                           RF_RD2_ADD_2_port, CK => Clk, Q => n_1082, QN => 
                           n1153);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx21x : DFF_X1 port map( D => n1558, CK 
                           => Clk, Q => RF_RD2_ADD_1_port, QN => n1377);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx1x : DFF_X1 port map( D => 
                           RF_RD2_ADD_1_port, CK => Clk, Q => n1883, QN => 
                           n1155);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx20x : DFF_X1 port map( D => n1559, CK 
                           => Clk, Q => RF_RD2_ADD_0_port, QN => n1376);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx0x : DFF_X1 port map( D => 
                           RF_RD2_ADD_0_port, CK => Clk, Q => n_1083, QN => 
                           n1152);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx19x : DFF_X1 port map( D => n1560, CK 
                           => Clk, Q => RF_RD1_ADD_4_port, QN => n1375);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx4x : DFF_X1 port map( D => 
                           RF_RD1_ADD_4_port, CK => Clk, Q => n1893, QN => 
                           n1164);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx18x : DFF_X1 port map( D => n1561, CK 
                           => Clk, Q => RF_RD1_ADD_3_port, QN => n1374);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx3x : DFF_X1 port map( D => 
                           RF_RD1_ADD_3_port, CK => Clk, Q => n1894, QN => 
                           n1165);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx17x : DFF_X1 port map( D => n1562, CK 
                           => Clk, Q => RF_RD1_ADD_2_port, QN => n1373);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx16x : DFF_X1 port map( D => n1563, CK 
                           => Clk, Q => RF_RD1_ADD_1_port, QN => n1372);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx15x : DFF_X1 port map( D => n1564, CK 
                           => Clk, Q => RF_RD1_ADD_0_port, QN => n1371);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx14x : DFF_X1 port map( D => n1565, CK 
                           => Clk, Q => n1210, QN => n1637);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx13x : DFF_X1 port map( D => n1566, CK 
                           => Clk, Q => n_1084, QN => n1635);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx12x : DFF_X1 port map( D => n1567, CK 
                           => Clk, Q => n_1085, QN => n1634);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx11x : DFF_X1 port map( D => n1568, CK 
                           => Clk, Q => DATAPATH_IxINSTR_11_port, QN => n1370);
   DATAPATH_IxSecond_stxWRADD_d1_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_11_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, QN => n_1086);
   DATAPATH_IxSecond_stxWRADD_d2_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_4_port, QN => n1150);
   DATAPATH_IxSecond_stxWRADD_d3_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_4_port, CK => Clk, Q => 
                           n2365, QN => n1158);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx10x : DFF_X1 port map( D => n1569, CK 
                           => Clk, Q => DATAPATH_IxINSTR_10_port, QN => n1369);
   DATAPATH_IxSecond_stxWRADD_d1_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_10_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, QN => n_1087);
   DATAPATH_IxSecond_stxWRADD_d2_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_3_port, QN => n_1088);
   DATAPATH_IxSecond_stxWRADD_d3_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_3_port, CK => Clk, Q => 
                           RF_WR_ADD(3), QN => n1160);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx9x : DFF_X1 port map( D => n1570, CK =>
                           Clk, Q => DATAPATH_IxINSTR_9_port, QN => n1368);
   DATAPATH_IxSecond_stxWRADD_d1_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_9_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, QN => n_1089);
   DATAPATH_IxSecond_stxWRADD_d2_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_2_port, QN => n1147);
   DATAPATH_IxSecond_stxWRADD_d3_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_2_port, CK => Clk, Q => 
                           RF_WR_ADD(2), QN => n1146);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx8x : DFF_X1 port map( D => n1571, CK =>
                           Clk, Q => DATAPATH_IxINSTR_8_port, QN => n1367);
   DATAPATH_IxSecond_stxWRADD_d1_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_8_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, QN => n_1090);
   DATAPATH_IxSecond_stxWRADD_d2_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_1_port, QN => n1148);
   DATAPATH_IxSecond_stxWRADD_d3_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_1_port, CK => Clk, Q => 
                           RF_WR_ADD(1), QN => n1159);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx7x : DFF_X1 port map( D => n1572, CK =>
                           Clk, Q => DATAPATH_IxINSTR_7_port, QN => n1366);
   DATAPATH_IxSecond_stxWRADD_d1_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_7_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, QN => n_1091);
   DATAPATH_IxSecond_stxWRADD_d2_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_0_port, QN => n1151);
   DATAPATH_IxSecond_stxWRADD_d3_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_0_port, CK => Clk, Q => 
                           RF_WR_ADD(0), QN => n1145);
   CU_Ixcw2_i_regx14x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1991, Q => n_1092, QN => n1211);
   CU_Ixcw2_i_regx12x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1991, Q => CU_Ixcw2_i_12_port, QN => n_1093);
   CU_Ixcw2_i_regx13x : DFFR_X1 port map( D => CU_Ixcw1_14_port, CK => Clk, RN 
                           => n1991, Q => n_1094, QN => n1212);
   CU_Ixcw2_i_regx8x : DFFR_X1 port map( D => CU_Ixcw1_8_port, CK => Clk, RN =>
                           n1991, Q => n_1095, QN => n1206);
   CU_Ixcw2_i_regx7x : DFFR_X1 port map( D => CU_Ixcw1_7_port, CK => Clk, RN =>
                           n1992, Q => n_1096, QN => n1207);
   CU_Ixcw2_i_regx5x : DFFR_X1 port map( D => CU_Ixcw1_5_port, CK => Clk, RN =>
                           n1992, Q => n_1097, QN => n1203);
   CU_Ixcw3_regx5x : DFFR_X1 port map( D => CU_Ixcw2_5_port, CK => Clk, RN => 
                           n1992, Q => IMM_SEL_i, QN => n1693);
   CU_Ixcw2_i_regx4x : DFFR_X1 port map( D => CU_Ixcw1_4_port, CK => Clk, RN =>
                           n1992, Q => n_1098, QN => n1202);
   CU_Ixcw3_regx4x : DFFR_X1 port map( D => CU_Ixcw2_4_port, CK => Clk, RN => 
                           n1992, Q => BRANCH_EN_i, QN => n_1099);
   CU_Ixcw2_i_regx9x : DFFR_X1 port map( D => CU_Ixcw1_9_port, CK => Clk, RN =>
                           n1992, Q => n_1100, QN => n1205);
   CU_Ixcw2_i_regx3x : DFFR_X1 port map( D => CU_Ixcw1_9_port, CK => Clk, RN =>
                           n1992, Q => n_1101, QN => n1201);
   CU_Ixcw3_regx3x : DFFR_X1 port map( D => CU_Ixcw2_3_port, CK => Clk, RN => 
                           n1992, Q => CU_Ixcw3_3_port, QN => n_1102);
   CU_Ixcw4_regx3x : DFFR_X1 port map( D => CU_Ixcw3_3_port, CK => Clk, RN => 
                           n1992, Q => DRAM_WE, QN => n_1103);
   CU_Ixcw2_i_regx2x : DFFR_X1 port map( D => CU_Ixcw1_2_port, CK => Clk, RN =>
                           n1992, Q => n_1104, QN => n1200);
   CU_Ixcw3_regx2x : DFFR_X1 port map( D => CU_Ixcw2_2_port, CK => Clk, RN => 
                           n1992, Q => CU_Ixcw3_2_port, QN => n_1105);
   CU_Ixcw4_regx2x : DFFR_X1 port map( D => CU_Ixcw3_2_port, CK => Clk, RN => 
                           n1991, Q => DRAM_RE, QN => n_1106);
   CU_Ixcw2_i_regx1x : DFFR_X1 port map( D => CU_Ixcw1_1_port, CK => Clk, RN =>
                           n1992, Q => n_1107, QN => n1199);
   CU_Ixcw3_regx1x : DFFR_X1 port map( D => CU_Ixcw2_1_port, CK => Clk, RN => 
                           n1992, Q => CU_Ixcw3_1_port, QN => n_1108);
   CU_Ixcw4_regx1x : DFFR_X1 port map( D => CU_Ixcw3_1_port, CK => Clk, RN => 
                           n1991, Q => WB_MUX_SEL_MEM_i, QN => n1334);
   CU_Ixcw2_i_regx6x : DFFR_X1 port map( D => CU_Ixcw1_6_port, CK => Clk, RN =>
                           n1992, Q => n_1109, QN => n1204);
   CU_Ixcw3_regx6x : DFFR_X1 port map( D => CU_Ixcw2_6_port, CK => Clk, RN => 
                           n1992, Q => PC_SEL_i, QN => n_1110);
   CU_Ixcw2_i_regx11x : DFFR_X1 port map( D => CU_Ixcw1_6_port, CK => Clk, RN 
                           => n1992, Q => CU_Ixcw2_i_11_port, QN => n_1111);
   CU_Ixcw2_i_regx10x : DFFR_X1 port map( D => CU_Ixcw1_10_port, CK => Clk, RN 
                           => n1992, Q => CU_Ixcw2_i_10_port, QN => n_1112);
   DATAPATH_IxSecond_stxIMM_out_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_4_port, CK => Clk,
                           Q => n_1113, QN => n1192);
   DATAPATH_IxSecond_stxIMM_out_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_3_port, CK => Clk,
                           Q => n_1114, QN => n1196);
   DATAPATH_IxSecond_stxIMM_out_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_2_port, CK => Clk,
                           Q => n_1115, QN => n1195);
   DATAPATH_IxSecond_stxIMM_out_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_1_port, CK => Clk,
                           Q => n_1116, QN => n1194);
   DATAPATH_IxSecond_stxIMM_out_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_31_port, CK => Clk
                           , Q => n_1117, QN => n1170);
   DATAPATH_IxSecond_stxIMM_out_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_30_port, CK => Clk
                           , Q => n_1118, QN => n1169);
   DATAPATH_IxSecond_stxIMM_out_regx29x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_29_port, CK => Clk
                           , Q => n_1119, QN => n1157);
   DATAPATH_IxSecond_stxIMM_out_regx28x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_28_port, CK => Clk
                           , Q => n_1120, QN => n1166);
   DATAPATH_IxSecond_stxIMM_out_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_27_port, CK => Clk
                           , Q => n_1121, QN => n1167);
   DATAPATH_IxSecond_stxIMM_out_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_26_port, CK => Clk
                           , Q => n_1122, QN => n1168);
   DATAPATH_IxSecond_stxIMM_out_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_25_port, CK => Clk
                           , Q => n_1123, QN => n1171);
   DATAPATH_IxSecond_stxIMM_out_regx24x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_24_port, CK => Clk
                           , Q => n_1124, QN => n1172);
   DATAPATH_IxSecond_stxIMM_out_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_23_port, CK => Clk
                           , Q => n_1125, QN => n1174);
   DATAPATH_IxSecond_stxIMM_out_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_22_port, CK => Clk
                           , Q => n_1126, QN => n1179);
   DATAPATH_IxSecond_stxIMM_out_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_21_port, CK => Clk
                           , Q => n_1127, QN => n1173);
   DATAPATH_IxSecond_stxIMM_out_regx20x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_20_port, CK => Clk
                           , Q => n_1128, QN => n1178);
   DATAPATH_IxSecond_stxIMM_out_regx19x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_19_port, CK => Clk
                           , Q => n_1129, QN => n1177);
   DATAPATH_IxSecond_stxIMM_out_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_18_port, CK => Clk
                           , Q => n_1130, QN => n1175);
   DATAPATH_IxSecond_stxIMM_out_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_17_port, CK => Clk
                           , Q => n_1131, QN => n1176);
   DATAPATH_IxSecond_stxIMM_out_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_16_port, CK => Clk
                           , Q => n_1132, QN => n1180);
   DATAPATH_IxSecond_stxIMM_out_regx15x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_15_port, CK => Clk
                           , Q => n_1133, QN => n1181);
   DATAPATH_IxSecond_stxIMM_out_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_14_port, CK => Clk
                           , Q => n_1134, QN => n1183);
   DATAPATH_IxSecond_stxIMM_out_regx13x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_13_port, CK => Clk
                           , Q => n_1135, QN => n1188);
   DATAPATH_IxSecond_stxIMM_out_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_12_port, CK => Clk
                           , Q => n_1136, QN => n1182);
   DATAPATH_IxSecond_stxIMM_out_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stximm_extended_0_port, CK => Clk,
                           Q => n_1137, QN => n1193);
   CU_Ixcw2_i_regx0x : DFFR_X1 port map( D => CU_Ixcw1_0_port, CK => Clk, RN =>
                           n1992, Q => n_1138, QN => n1198);
   CU_Ixcw3_regx0x : DFFR_X1 port map( D => CU_Ixcw2_0_port, CK => Clk, RN => 
                           n1992, Q => CU_Ixcw3_0_port, QN => n_1139);
   CU_Ixcw4_regx0x : DFFR_X1 port map( D => CU_Ixcw3_0_port, CK => Clk, RN => 
                           n1992, Q => RF_WE_MEM_i, QN => n1333);
   CU_Ixcw5_regx0x : DFFR_X1 port map( D => RF_WE_MEM_i, CK => Clk, RN => n1992
                           , Q => RF_WR_EN, QN => n1299);
   DATAPATH_IxFirst_stxPC_regx1x : DFF_X1 port map( D => n1546, CK => Clk, Q =>
                           DATAPATH_IxPC4_1_port, QN => n1388);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx1x : DFF_X1 port map( D => n1513, CK =>
                           Clk, Q => n1592, QN => n1339);
   DATAPATH_IxSecond_stxPC_out_regx1x : DFF_X1 port map( D => n1512, CK => Clk,
                           Q => n_1140, QN => n1610);
   DATAPATH_IxSecond_stxBR_target_regx1x : DFF_X1 port map( D => n2090, CK => 
                           Clk, Q => n_1141, QN => n1214);
   DATAPATH_IxFirst_stxPC_regx0x : DFF_X1 port map( D => n1547, CK => Clk, Q =>
                           DATAPATH_IxPC4_0_port, QN => n1387);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx0x : DFF_X1 port map( D => n1515, CK =>
                           Clk, Q => DATAPATH_IxSecond_stxjump_target_0_port, 
                           QN => n1338);
   DATAPATH_IxSecond_stxBR_target_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_0_port, CK => Clk, 
                           Q => n_1142, QN => n1213);
   DATAPATH_IxSecond_stxPC_out_regx0x : DFF_X1 port map( D => n1514, CK => Clk,
                           Q => n_1143, QN => n1625);
   DATAPATH_IxFirst_stxPC_regx2x : DFF_X1 port map( D => n1545, CK => Clk, Q =>
                           IRAM_ADD_2_port, QN => n1389);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx2x : DFF_X1 port map( D => n1511, CK =>
                           Clk, Q => n1241, QN => n1591);
   DATAPATH_IxSecond_stxPC_out_regx2x : DFF_X1 port map( D => n1510, CK => Clk,
                           Q => n_1144, QN => n1621);
   DATAPATH_IxSecond_stxBR_target_regx2x : DFF_X1 port map( D => n1296, CK => 
                           Clk, Q => DATAPATH_IxSecond_stxBR_target_2_port, QN 
                           => n_1145);
   DATAPATH_IxFirst_stxPC_regx3x : DFF_X1 port map( D => n1544, CK => Clk, Q =>
                           IRAM_ADD_3_port, QN => n1390);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx3x : DFF_X1 port map( D => n1509, CK =>
                           Clk, Q => n1782, QN => n1340);
   DATAPATH_IxSecond_stxPC_out_regx3x : DFF_X1 port map( D => n1508, CK => Clk,
                           Q => n_1146, QN => n1619);
   DATAPATH_IxSecond_stxBR_target_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_3_port, CK => Clk, 
                           Q => n_1147, QN => n1215);
   DATAPATH_IxFirst_stxPC_regx4x : DFF_X1 port map( D => n1543, CK => Clk, Q =>
                           IRAM_ADD_4_port, QN => n1391);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx4x : DFF_X1 port map( D => n1507, CK =>
                           Clk, Q => n1244, QN => n1645);
   DATAPATH_IxSecond_stxPC_out_regx4x : DFF_X1 port map( D => n1506, CK => Clk,
                           Q => n_1148, QN => n1598);
   DATAPATH_IxSecond_stxBR_target_regx4x : DFF_X1 port map( D => n2085, CK => 
                           Clk, Q => n_1149, QN => n1216);
   DATAPATH_IxFirst_stxPC_regx5x : DFF_X1 port map( D => n1542, CK => Clk, Q =>
                           IRAM_ADD_5_port, QN => n1392);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx5x : DFF_X1 port map( D => n1505, CK =>
                           Clk, Q => n_1150, QN => n1341);
   DATAPATH_IxSecond_stxBR_target_regx5x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_5_port, CK => Clk, 
                           Q => n_1151, QN => n1217);
   DATAPATH_IxSecond_stxPC_out_regx5x : DFF_X1 port map( D => n1504, CK => Clk,
                           Q => n_1152, QN => n1609);
   DATAPATH_IxFirst_stxPC_regx6x : DFF_X1 port map( D => n1541, CK => Clk, Q =>
                           IRAM_ADD_6_port, QN => n1393);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx6x : DFF_X1 port map( D => n1503, CK =>
                           Clk, Q => n_1153, QN => n1342);
   DATAPATH_IxSecond_stxBR_target_regx6x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_6_port, CK => Clk, 
                           Q => DATAPATH_IxSecond_stxBR_target_6_port, QN => 
                           n_1154);
   DATAPATH_IxSecond_stxPC_out_regx6x : DFF_X1 port map( D => n1502, CK => Clk,
                           Q => n_1155, QN => n1620);
   DATAPATH_IxFirst_stxPC_regx7x : DFF_X1 port map( D => n1540, CK => Clk, Q =>
                           IRAM_ADD_7_port, QN => n1394);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx7x : DFF_X1 port map( D => n1501, CK =>
                           Clk, Q => n1248, QN => n1636);
   DATAPATH_IxSecond_stxBR_target_regx7x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_7_port, CK => Clk, 
                           Q => n_1156, QN => n1218);
   DATAPATH_IxSecond_stxPC_out_regx7x : DFF_X1 port map( D => n1500, CK => Clk,
                           Q => n_1157, QN => n1599);
   DATAPATH_IxFirst_stxPC_regx8x : DFF_X1 port map( D => n1539, CK => Clk, Q =>
                           IRAM_ADD_8_port, QN => n1395);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx8x : DFF_X1 port map( D => n1499, CK =>
                           Clk, Q => n_1158, QN => n1343);
   DATAPATH_IxSecond_stxPC_out_regx8x : DFF_X1 port map( D => n1498, CK => Clk,
                           Q => n_1159, QN => n1594);
   DATAPATH_IxSecond_stxBR_target_regx8x : DFF_X1 port map( D => n1291, CK => 
                           Clk, Q => DATAPATH_IxSecond_stxBR_target_8_port, QN 
                           => n_1160);
   DATAPATH_IxFirst_stxPC_regx9x : DFF_X1 port map( D => n1538, CK => Clk, Q =>
                           IRAM_ADD_9_port, QN => n1396);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx9x : DFF_X1 port map( D => n1497, CK =>
                           Clk, Q => n_1161, QN => n1344);
   DATAPATH_IxSecond_stxPC_out_regx9x : DFF_X1 port map( D => n1496, CK => Clk,
                           Q => n_1162, QN => n1606);
   DATAPATH_IxSecond_stxBR_target_regx9x : DFF_X1 port map( D => n2082, CK => 
                           Clk, Q => n_1163, QN => n1219);
   DATAPATH_IxFirst_stxPC_regx10x : DFF_X1 port map( D => n1537, CK => Clk, Q 
                           => IRAM_ADD_10_port, QN => n1397);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx10x : DFF_X1 port map( D => n1495, CK 
                           => Clk, Q => n_1164, QN => n1345);
   DATAPATH_IxSecond_stxPC_out_regx10x : DFF_X1 port map( D => n1494, CK => Clk
                           , Q => n_1165, QN => n1629);
   DATAPATH_IxSecond_stxBR_target_regx10x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_10_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_10_port, QN => 
                           n_1166);
   DATAPATH_IxFirst_stxPC_regx11x : DFF_X1 port map( D => n1536, CK => Clk, Q 
                           => IRAM_ADD_11_port, QN => n1398);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx11x : DFF_X1 port map( D => n1493, CK 
                           => Clk, Q => n_1167, QN => n1346);
   DATAPATH_IxSecond_stxBR_target_regx11x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_11_port, CK => Clk,
                           Q => n_1168, QN => n1220);
   DATAPATH_IxSecond_stxPC_out_regx11x : DFF_X1 port map( D => n1492, CK => Clk
                           , Q => n_1169, QN => n1626);
   DATAPATH_IxFirst_stxPC_regx12x : DFF_X1 port map( D => n1535, CK => Clk, Q 
                           => IRAM_ADD_12_port, QN => n1399);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx12x : DFF_X1 port map( D => n1491, CK 
                           => Clk, Q => n_1170, QN => n1347);
   DATAPATH_IxSecond_stxPC_out_regx12x : DFF_X1 port map( D => n1490, CK => Clk
                           , Q => n_1171, QN => n1615);
   DATAPATH_IxSecond_stxBR_target_regx13x : DFF_X1 port map( D => n2068, CK => 
                           Clk, Q => n_1172, QN => n1221);
   DATAPATH_IxFirst_stxPC_regx13x : DFF_X1 port map( D => n1534, CK => Clk, Q 
                           => IRAM_ADD_13_port, QN => n1400);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx13x : DFF_X1 port map( D => n1489, CK 
                           => Clk, Q => n_1173, QN => n1348);
   DATAPATH_IxSecond_stxPC_out_regx13x : DFF_X1 port map( D => n1488, CK => Clk
                           , Q => n_1174, QN => n1630);
   DATAPATH_IxFirst_stxPC_regx14x : DFF_X1 port map( D => n1533, CK => Clk, Q 
                           => IRAM_ADD_14_port, QN => n1401);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx14x : DFF_X1 port map( D => n1487, CK 
                           => Clk, Q => n1641, QN => n1349);
   DATAPATH_IxSecond_stxPC_out_regx14x : DFF_X1 port map( D => n1486, CK => Clk
                           , Q => n_1175, QN => n1596);
   DATAPATH_IxSecond_stxBR_target_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_14_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_14_port, QN => 
                           n_1176);
   DATAPATH_IxFirst_stxPC_regx15x : DFF_X1 port map( D => n1532, CK => Clk, Q 
                           => IRAM_ADD_15_port, QN => n1402);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx15x : DFF_X1 port map( D => n1485, CK 
                           => Clk, Q => n1257, QN => n1707);
   DATAPATH_IxSecond_stxPC_out_regx15x : DFF_X1 port map( D => n1484, CK => Clk
                           , Q => n_1177, QN => n1593);
   DATAPATH_IxSecond_stxBR_target_regx15x : DFF_X1 port map( D => n2066, CK => 
                           Clk, Q => n_1178, QN => n1222);
   DATAPATH_IxSecond_stxBR_target_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_12_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_12_port, QN => 
                           n_1179);
   DATAPATH_IxSecond_stxBR_target_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_16_port, CK => Clk,
                           Q => n_1180, QN => n1223);
   DATAPATH_IxFirst_stxPC_regx16x : DFF_X1 port map( D => n1531, CK => Clk, Q 
                           => IRAM_ADD_16_port, QN => n1403);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx16x : DFF_X1 port map( D => n1483, CK 
                           => Clk, Q => n_1181, QN => n1350);
   DATAPATH_IxSecond_stxPC_out_regx16x : DFF_X1 port map( D => n1482, CK => Clk
                           , Q => n_1182, QN => n1597);
   DATAPATH_IxSecond_stxBR_target_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_17_port, CK => Clk,
                           Q => n_1183, QN => n1224);
   DATAPATH_IxFirst_stxPC_regx17x : DFF_X1 port map( D => n1530, CK => Clk, Q 
                           => IRAM_ADD_17_port, QN => n1404);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx17x : DFF_X1 port map( D => n1481, CK 
                           => Clk, Q => n_1184, QN => n1351);
   DATAPATH_IxSecond_stxPC_out_regx17x : DFF_X1 port map( D => n1480, CK => Clk
                           , Q => n_1185, QN => n1604);
   DATAPATH_IxSecond_stxBR_target_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_18_port, CK => Clk,
                           Q => DATAPATH_IxSecond_stxBR_target_18_port, QN => 
                           n_1186);
   DATAPATH_IxFirst_stxPC_regx18x : DFF_X1 port map( D => n1529, CK => Clk, Q 
                           => IRAM_ADD_18_port, QN => n1405);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx18x : DFF_X1 port map( D => n1479, CK 
                           => Clk, Q => n_1187, QN => n1352);
   DATAPATH_IxSecond_stxPC_out_regx18x : DFF_X1 port map( D => n1478, CK => Clk
                           , Q => n_1188, QN => n1611);
   DATAPATH_IxFirst_stxPC_regx19x : DFF_X1 port map( D => n1528, CK => Clk, Q 
                           => IRAM_ADD_19_port, QN => n1406);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx19x : DFF_X1 port map( D => n1477, CK 
                           => Clk, Q => n_1189, QN => n1353);
   DATAPATH_IxSecond_stxBR_target_regx19x : DFF_X1 port map( D => n2050, CK => 
                           Clk, Q => n_1190, QN => n1225);
   DATAPATH_IxSecond_stxPC_out_regx19x : DFF_X1 port map( D => n1476, CK => Clk
                           , Q => n_1191, QN => n1600);
   DATAPATH_IxFirst_stxPC_regx20x : DFF_X1 port map( D => n1527, CK => Clk, Q 
                           => IRAM_ADD_20_port, QN => n1407);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx20x : DFF_X1 port map( D => n1475, CK 
                           => Clk, Q => n_1192, QN => n1354);
   DATAPATH_IxSecond_stxPC_out_regx20x : DFF_X1 port map( D => n1474, CK => Clk
                           , Q => n_1193, QN => n1612);
   DATAPATH_IxSecond_stxBR_target_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_21_port, CK => Clk,
                           Q => n_1194, QN => n1227);
   DATAPATH_IxFirst_stxPC_regx21x : DFF_X1 port map( D => n1526, CK => Clk, Q 
                           => IRAM_ADD_21_port, QN => n1408);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx21x : DFF_X1 port map( D => n1473, CK 
                           => Clk, Q => n_1195, QN => n1355);
   DATAPATH_IxSecond_stxPC_out_regx21x : DFF_X1 port map( D => n1472, CK => Clk
                           , Q => n_1196, QN => n1618);
   DATAPATH_IxSecond_stxBR_target_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_22_port, CK => Clk,
                           Q => n_1197, QN => n1228);
   DATAPATH_IxFirst_stxPC_regx22x : DFF_X1 port map( D => n1525, CK => Clk, Q 
                           => IRAM_ADD_22_port, QN => n1409);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx22x : DFF_X1 port map( D => n1471, CK 
                           => Clk, Q => n1639, QN => n1356);
   DATAPATH_IxSecond_stxPC_out_regx22x : DFF_X1 port map( D => n1470, CK => Clk
                           , Q => n_1198, QN => n1614);
   DATAPATH_IxSecond_stxBR_target_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_23_port, CK => Clk,
                           Q => n_1199, QN => n1229);
   DATAPATH_IxFirst_stxPC_regx23x : DFF_X1 port map( D => n1524, CK => Clk, Q 
                           => IRAM_ADD_23_port, QN => n1410);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx23x : DFF_X1 port map( D => n1469, CK 
                           => Clk, Q => n_1200, QN => n1357);
   DATAPATH_IxSecond_stxPC_out_regx23x : DFF_X1 port map( D => n1468, CK => Clk
                           , Q => n_1201, QN => n1617);
   DATAPATH_IxSecond_stxBR_target_regx20x : DFF_X1 port map( D => n1292, CK => 
                           Clk, Q => n_1202, QN => n1226);
   DATAPATH_IxSecond_stxBR_target_regx24x : DFF_X1 port map( D => n2054, CK => 
                           Clk, Q => n_1203, QN => n1230);
   DATAPATH_IxFirst_stxPC_regx24x : DFF_X1 port map( D => n1523, CK => Clk, Q 
                           => IRAM_ADD_24_port, QN => n1411);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx24x : DFF_X1 port map( D => n1467, CK 
                           => Clk, Q => n_1204, QN => n1358);
   DATAPATH_IxSecond_stxPC_out_regx24x : DFF_X1 port map( D => n1466, CK => Clk
                           , Q => n_1205, QN => n1595);
   DATAPATH_IxSecond_stxBR_target_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_25_port, CK => Clk,
                           Q => n_1206, QN => n1231);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx25x : DFF_X1 port map( D => n1465, CK 
                           => Clk, Q => n_1207, QN => n1359);
   DATAPATH_IxSecond_stxPC_out_regx25x : DFF_X1 port map( D => n1464, CK => Clk
                           , Q => n_1208, QN => n1613);
   DATAPATH_IxFirst_stxPC_regx26x : DFF_X1 port map( D => n1521, CK => Clk, Q 
                           => IRAM_ADD_26_port, QN => n1413);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx26x : DFF_X1 port map( D => n1463, CK 
                           => Clk, Q => n1640, QN => n1360);
   DATAPATH_IxSecond_stxPC_out_regx26x : DFF_X1 port map( D => n1462, CK => Clk
                           , Q => n_1209, QN => n1627);
   DATAPATH_IxSecond_stxBR_target_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_26_port, CK => Clk,
                           Q => n_1210, QN => n1232);
   DATAPATH_IxFirst_stxPC_regx27x : DFF_X1 port map( D => n1520, CK => Clk, Q 
                           => IRAM_ADD_27_port, QN => n1414);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx27x : DFF_X1 port map( D => n1461, CK 
                           => Clk, Q => n_1211, QN => n1361);
   DATAPATH_IxSecond_stxBR_target_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_27_port, CK => Clk,
                           Q => n_1212, QN => n1233);
   DATAPATH_IxSecond_stxPC_out_regx27x : DFF_X1 port map( D => n1460, CK => Clk
                           , Q => n_1213, QN => n1628);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx28x : DFF_X1 port map( D => n1459, CK 
                           => Clk, Q => n1690, QN => n1362);
   DATAPATH_IxSecond_stxPC_out_regx28x : DFF_X1 port map( D => n1458, CK => Clk
                           , Q => n_1214, QN => n1608);
   DATAPATH_IxSecond_stxBR_target_regx29x : DFF_X1 port map( D => n2061, CK => 
                           Clk, Q => n_1215, QN => n1235);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx29x : DFF_X1 port map( D => n1457, CK 
                           => Clk, Q => n_1216, QN => n1363);
   DATAPATH_IxSecond_stxPC_out_regx29x : DFF_X1 port map( D => n1456, CK => Clk
                           , Q => n_1217, QN => n1607);
   DATAPATH_IxSecond_stxBR_target_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_30_port, CK => Clk,
                           Q => n_1218, QN => n1236);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx30x : DFF_X1 port map( D => n1455, CK 
                           => Clk, Q => n1638, QN => n1364);
   DATAPATH_IxSecond_stxPC_out_regx30x : DFF_X1 port map( D => n1454, CK => Clk
                           , Q => n_1219, QN => n1616);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_1_port, CK => Clk, Q 
                           => DRAM_ADD_1_port, QN => n1420);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx1x : DFF_X1 port map( D => 
                           DRAM_ADD_1_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_1_port, QN => n_1220);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_2_port, CK => Clk, Q 
                           => DRAM_ADD_2_port, QN => n1421);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx2x : DFF_X1 port map( D => 
                           DRAM_ADD_2_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_2_port, QN => n_1221);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_3_port, CK => Clk, Q 
                           => DRAM_ADD_3_port, QN => n1422);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx3x : DFF_X1 port map( D => 
                           DRAM_ADD_3_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_3_port, QN => n_1222);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_4_port, CK => Clk, Q 
                           => DRAM_ADD_4_port, QN => n1423);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx4x : DFF_X1 port map( D => 
                           DRAM_ADD_4_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_4_port, QN => n_1223);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx5x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_5_port, CK => Clk, Q 
                           => DRAM_ADD_5_port, QN => n1424);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx5x : DFF_X1 port map( D => 
                           DRAM_ADD_5_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_5_port, QN => n_1224);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx6x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_6_port, CK => Clk, Q 
                           => DRAM_ADD_6_port, QN => n1425);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx6x : DFF_X1 port map( D => 
                           DRAM_ADD_6_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_6_port, QN => n_1225);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx7x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_7_port, CK => Clk, Q 
                           => DRAM_ADD_7_port, QN => n1426);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx7x : DFF_X1 port map( D => 
                           DRAM_ADD_7_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_7_port, QN => n_1226);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx8x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_8_port, CK => Clk, Q 
                           => DRAM_ADD_8_port, QN => n1427);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx8x : DFF_X1 port map( D => 
                           DRAM_ADD_8_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_8_port, QN => n_1227);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx9x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_9_port, CK => Clk, Q 
                           => DRAM_ADD_9_port, QN => n1428);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx9x : DFF_X1 port map( D => 
                           DRAM_ADD_9_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_9_port, QN => n_1228);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx11x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_11_port, CK => Clk, Q 
                           => DRAM_ADD_11_port, QN => n1430);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx11x : DFF_X1 port map( D => 
                           DRAM_ADD_11_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_11_port, QN => n_1229);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_12_port, CK => Clk, Q 
                           => DRAM_ADD_12_port, QN => n1431);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx12x : DFF_X1 port map( D => 
                           DRAM_ADD_12_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_12_port, QN => n_1230);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx13x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_13_port, CK => Clk, Q 
                           => DRAM_ADD_13_port, QN => n1432);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx13x : DFF_X1 port map( D => 
                           DRAM_ADD_13_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_13_port, QN => n_1231);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_14_port, CK => Clk, Q 
                           => DRAM_ADD_14_port, QN => n1433);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx14x : DFF_X1 port map( D => 
                           DRAM_ADD_14_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_14_port, QN => n_1232);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx15x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_15_port, CK => Clk, Q 
                           => DRAM_ADD_15_port, QN => n1434);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx15x : DFF_X1 port map( D => 
                           DRAM_ADD_15_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_15_port, QN => n_1233);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx19x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_19_port, CK => Clk, Q 
                           => DRAM_ADD_19_port, QN => n1438);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx19x : DFF_X1 port map( D => 
                           DRAM_ADD_19_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_19_port, QN => n_1234);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx20x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_20_port, CK => Clk, Q 
                           => DRAM_ADD_20_port, QN => n1439);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx20x : DFF_X1 port map( D => 
                           DRAM_ADD_20_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_20_port, QN => n_1235);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_21_port, CK => Clk, Q 
                           => DRAM_ADD_21_port, QN => n1440);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx21x : DFF_X1 port map( D => 
                           DRAM_ADD_21_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_21_port, QN => n_1236);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_22_port, CK => Clk, Q 
                           => DRAM_ADD_22_port, QN => n1441);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx22x : DFF_X1 port map( D => 
                           DRAM_ADD_22_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_22_port, QN => n_1237);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_23_port, CK => Clk, Q 
                           => DRAM_ADD_23_port, QN => n1442);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx23x : DFF_X1 port map( D => 
                           DRAM_ADD_23_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_23_port, QN => n_1238);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx24x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_24_port, CK => Clk, Q 
                           => DRAM_ADD_24_port, QN => n1443);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx24x : DFF_X1 port map( D => 
                           DRAM_ADD_24_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_24_port, QN => n_1239);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_27_port, CK => Clk, Q 
                           => DRAM_ADD_27_port, QN => n1446);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx27x : DFF_X1 port map( D => 
                           DRAM_ADD_27_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_27_port, QN => n_1240);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx28x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_28_port, CK => Clk, Q 
                           => DRAM_ADD_28_port, QN => n1447);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx28x : DFF_X1 port map( D => 
                           DRAM_ADD_28_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_28_port, QN => n_1241);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx29x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_29_port, CK => Clk, Q 
                           => DRAM_ADD_29_port, QN => n1448);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx29x : DFF_X1 port map( D => 
                           DRAM_ADD_29_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_29_port, QN => n_1242);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_30_port, CK => Clk, Q 
                           => DRAM_ADD_30_port, QN => n1449);
   DATAPATH_IxFourth_stxALU_FORWARD_out_regx30x : DFF_X1 port map( D => 
                           DRAM_ADD_30_port, CK => Clk, Q => 
                           DATAPATH_IxALUOUT_Data1_30_port, QN => n_1243);
   DATAPATH_IxSecond_stxBR_target_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxjump_target_31_port, CK => Clk,
                           Q => n_1244, QN => n1237);
   DATAPATH_IxFirst_stxLATCH_PC_out_regx31x : DFF_X1 port map( D => n1453, CK 
                           => Clk, Q => n_1245, QN => n1365);
   DATAPATH_IxSecond_stxPC_out_regx31x : DFF_X1 port map( D => n1452, CK => Clk
                           , Q => n_1246, QN => n1622);
   DATAPATH_IxSecond_stxBR_target_regx28x : DFF_X1 port map( D => n2058, CK => 
                           Clk, Q => n_1247, QN => n1234);
   U5 : NAND3_X1 port map( A1 => n22, A2 => n23, A3 => n2002, ZN => n1287);
   U10 : NAND3_X1 port map( A1 => n32, A2 => n33, A3 => n2003, ZN => n1288);
   U13 : NAND3_X1 port map( A1 => n33, A2 => n23, A3 => n36, ZN => n1289);
   U19 : NAND3_X1 port map( A1 => IRAM_DOUT(14), A2 => IRAM_DOUT(12), A3 => n43
                           , ZN => n32);
   U22 : NAND3_X1 port map( A1 => IRAM_DOUT(5), A2 => n28, A3 => IRAM_DOUT(2), 
                           ZN => n33);
   U115 : NAND3_X1 port map( A1 => IRAM_ADD_28_port, A2 => IRAM_ADD_27_port, A3
                           => n118, ZN => n110);
   U153 : XOR2_X1 port map( A => n2057, B => n152, Z => n46);
   U165 : XOR2_X1 port map( A => n1409, B => n164, Z => n162);
   U182 : XOR2_X1 port map( A => n180, B => n1859, Z => n1292);
   U280 : XOR2_X1 port map( A => n268, B => n269, Z => n48);
   U304 : NAND3_X1 port map( A1 => n2095, A2 => n165, A3 => n1992, ZN => n289);
   U387 : XOR2_X1 port map( A => n358, B => n359, Z => n356);
   U389 : XOR2_X1 port map( A => n363, B => n359, Z => n355);
   U397 : XOR2_X1 port map( A => n360, B => n375, Z => n374);
   U399 : XOR2_X1 port map( A => n364, B => n375, Z => n373);
   U404 : XOR2_X1 port map( A => n386, B => n387, Z => n383);
   U416 : XOR2_X1 port map( A => n403, B => n404, Z => n402);
   U430 : XOR2_X1 port map( A => n432, B => n433, Z => n431);
   U431 : XOR2_X1 port map( A => n434, B => n433, Z => n428);
   U457 : XOR2_X1 port map( A => n474, B => n475, Z => n473);
   U459 : XOR2_X1 port map( A => n479, B => n475, Z => n470);
   U467 : XOR2_X1 port map( A => n476, B => n491, Z => n490);
   U469 : NAND3_X1 port map( A1 => n2104, A2 => n1785, A3 => n495, ZN => n493);
   U471 : XOR2_X1 port map( A => n480, B => n491, Z => n489);
   U477 : XOR2_X1 port map( A => n504, B => n505, Z => n501);
   U491 : XOR2_X1 port map( A => n523, B => n524, Z => n522);
   U493 : XOR2_X1 port map( A => n528, B => n524, Z => n519);
   U500 : XOR2_X1 port map( A => n525, B => n539, Z => n538);
   U502 : NAND3_X1 port map( A1 => n2108, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, A3 => n543, ZN 
                           => n541);
   U504 : XOR2_X1 port map( A => n529, B => n539, Z => n537);
   U510 : XOR2_X1 port map( A => n552, B => n553, Z => n549);
   U523 : XOR2_X1 port map( A => n442, B => n1743, Z => n567);
   U533 : XOR2_X1 port map( A => n581, B => n582, Z => n579);
   U535 : XOR2_X1 port map( A => n586, B => n582, Z => n578);
   U542 : XOR2_X1 port map( A => n583, B => n597, Z => n596);
   U545 : XOR2_X1 port map( A => n587, B => n597, Z => n595);
   U566 : XOR2_X1 port map( A => n629, B => n630, Z => n628);
   U568 : XOR2_X1 port map( A => n634, B => n630, Z => n625);
   U575 : XOR2_X1 port map( A => n631, B => n645, Z => n644);
   U577 : XOR2_X1 port map( A => n635, B => n645, Z => n643);
   U582 : XOR2_X1 port map( A => n656, B => n657, Z => n653);
   U594 : XOR2_X1 port map( A => n673, B => n674, Z => n672);
   U596 : XOR2_X1 port map( A => n678, B => n674, Z => n671);
   U603 : XOR2_X1 port map( A => n675, B => n689, Z => n688);
   U606 : XOR2_X1 port map( A => n679, B => n689, Z => n687);
   U608 : NAND3_X1 port map( A1 => n2119, A2 => n1809, A3 => n337, ZN => n693);
   U615 : NAND3_X1 port map( A1 => n1335, A2 => n1930, A3 => n1336, ZN => n418)
                           ;
   U625 : XOR2_X1 port map( A => n707, B => n420, Z => n706);
   U628 : XOR2_X1 port map( A => n420, B => n712, Z => n710);
   U695 : XOR2_X1 port map( A => n1921, B => n1580, Z => n657);
   U699 : XOR2_X1 port map( A => n1921, B => n2152, Z => n658);
   U710 : XOR2_X1 port map( A => n1921, B => n333, Z => n336);
   U725 : XOR2_X1 port map( A => n1921, B => n1985, Z => n388);
   U727 : XOR2_X1 port map( A => n1921, B => n1739, Z => n404);
   U750 : XOR2_X1 port map( A => n1921, B => n663, Z => n664);
   U767 : XOR2_X1 port map( A => n1921, B => n610, Z => n783);
   U783 : XOR2_X1 port map( A => n791, B => n792, Z => n237);
   U787 : XOR2_X1 port map( A => n798, B => n799, Z => n797);
   U789 : XOR2_X1 port map( A => n803, B => n799, Z => n795);
   U794 : XOR2_X1 port map( A => n800, B => n808, Z => n807);
   U796 : XOR2_X1 port map( A => n804, B => n808, Z => n806);
   U798 : XOR2_X1 port map( A => n812, B => n813, Z => 
                           DATAPATH_IxSecond_stxjump_target_5_port);
   U804 : XOR2_X1 port map( A => n821, B => n822, Z => n820);
   U806 : XOR2_X1 port map( A => n825, B => n822, Z => n818);
   U807 : XOR2_X1 port map( A => n1365, B => n1386, Z => n822);
   U811 : XOR2_X1 port map( A => n829, B => n824, Z => n828);
   U813 : XOR2_X1 port map( A => n826, B => n829, Z => n827);
   U834 : XOR2_X1 port map( A => n838, B => n843, Z => n847);
   U836 : XOR2_X1 port map( A => n845, B => n838, Z => n846);
   U856 : XOR2_X1 port map( A => n854, B => n860, Z => n864);
   U858 : XOR2_X1 port map( A => n862, B => n854, Z => n863);
   U872 : XOR2_X1 port map( A => n879, B => n869, Z => n182);
   U888 : XOR2_X1 port map( A => n898, B => n874, Z => 
                           DATAPATH_IxSecond_stxjump_target_17_port);
   U915 : XOR2_X1 port map( A => n905, B => n910, Z => n920);
   U917 : XOR2_X1 port map( A => n905, B => n917, Z => n918);
   U937 : XOR2_X1 port map( A => n1384, B => n1343, Z => n244);
   U946 : XOR2_X1 port map( A => n940, B => n930, Z => n939);
   U948 : XOR2_X1 port map( A => n944, B => n930, Z => n938);
   U955 : XOR2_X1 port map( A => n942, B => n931, Z => n948);
   U958 : XOR2_X1 port map( A => n946, B => n931, Z => n947);
   U963 : NAND3_X1 port map( A1 => n1343, A2 => n2196, A3 => n1384, ZN => n951)
                           ;
   U969 : XOR2_X1 port map( A => n1383, B => n1248, Z => n799);
   U999 : XOR2_X1 port map( A => n1382, B => n1342, Z => n808);
   U1192 : XOR2_X1 port map( A => n2134, B => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, Z => n463);
   U1341 : NAND3_X1 port map( A1 => n1930, A2 => n1605, A3 => n1335, ZN => n790
                           );
   U1353 : XOR2_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_1_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, Z => n565);
   U1377 : XOR2_X1 port map( A => n1160, B => n1165, Z => n1106);
   U1401 : XOR2_X1 port map( A => n1147, B => n1153, Z => n1124);
   U1422 : NAND3_X1 port map( A1 => n1134, A2 => n26, A3 => n1139, ZN => 
                           CU_IxN24);
   U310 : NOR3_X2 port map( A1 => n1993, A2 => n109, A3 => n165, ZN => n190);
   U978 : AND2_X2 port map( A1 => n1244, A2 => n956, ZN => n270);
   U1363 : OAI21_X2 port map( B1 => n1810, B2 => PC_SEL_i, A => n1092, ZN => 
                           n1088);
   DATAPATH_IxFirst_stxPC_regx30x : DFF_X1 port map( D => n1517, CK => Clk, Q 
                           => IRAM_ADD_30_port, QN => n1417);
   DATAPATH_IxFirst_stxPC_regx31x : DFF_X1 port map( D => n1516, CK => Clk, Q 
                           => IRAM_ADD_31_port, QN => n1418);
   DATAPATH_IxFirst_stxPC_regx28x : DFF_X1 port map( D => n1519, CK => Clk, Q 
                           => IRAM_ADD_28_port, QN => n1415);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_0_port, CK => Clk, Q 
                           => DRAM_ADD_0_port, QN => n1419);
   DATAPATH_IxFirst_stxPC_regx29x : DFF_X1 port map( D => n1518, CK => Clk, Q 
                           => IRAM_ADD_29_port, QN => n1416);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx2x : DFF_X1 port map( D => 
                           RF_RD1_ADD_2_port, CK => Clk, Q => n1895, QN => 
                           n1163);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx1x : DFF_X1 port map( D => 
                           RF_RD1_ADD_1_port, CK => Clk, Q => n1811, QN => 
                           n1877);
   DATAPATH_IxSecond_stxRF_ADD_RD1_EX_regx0x : DFF_X1 port map( D => 
                           RF_RD1_ADD_0_port, CK => Clk, Q => n1813, QN => 
                           n1878);
   DATAPATH_IxSecond_stxRF_ADD_RD2_EX_regx3x : DFF_X1 port map( D => 
                           RF_RD2_ADD_3_port, CK => Clk, Q => n1887, QN => 
                           n1156);
   DATAPATH_IxSecond_stxIMM_out_regx11x : DFF_X1 port map( D => n1688, CK => 
                           Clk, Q => n_1248, QN => n1187);
   DATAPATH_IxSecond_stxIMM_out_regx10x : DFF_X1 port map( D => n1687, CK => 
                           Clk, Q => n_1249, QN => n1186);
   DATAPATH_IxSecond_stxIMM_out_regx9x : DFF_X1 port map( D => n1686, CK => Clk
                           , Q => n_1250, QN => n1184);
   DATAPATH_IxSecond_stxIMM_out_regx8x : DFF_X1 port map( D => n1685, CK => Clk
                           , Q => n_1251, QN => n1185);
   DATAPATH_IxSecond_stxIMM_out_regx7x : DFF_X1 port map( D => n1684, CK => Clk
                           , Q => n_1252, QN => n1189);
   DATAPATH_IxSecond_stxIMM_out_regx6x : DFF_X1 port map( D => n1683, CK => Clk
                           , Q => n_1253, QN => n1190);
   DATAPATH_IxSecond_stxIMM_out_regx5x : DFF_X1 port map( D => n1682, CK => Clk
                           , Q => n_1254, QN => n1191);
   CU_Ixcw5_regx1x : DFFR_X1 port map( D => WB_MUX_SEL_MEM_i, CK => Clk, RN => 
                           n1992, Q => n1939, QN => n1590);
   DATAPATH_IxFirst_stxPC_regx25x : DFF_X1 port map( D => n1522, CK => Clk, Q 
                           => IRAM_ADD_25_port, QN => n1412);
   U1445 : XNOR2_X1 port map( A => n1711, B => n1573, ZN => n47);
   U1446 : XOR2_X1 port map( A => n1362, B => n1914, Z => n1573);
   U1447 : OAI221_X4 port map( B1 => n1871, B2 => n1599, C1 => n1426, C2 => 
                           n1823, A => n1064, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_7_port);
   U1448 : OAI221_X4 port map( B1 => n1871, B2 => n1610, C1 => n1420, C2 => 
                           n1823, A => n1086, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_1_port);
   U1449 : OAI221_X4 port map( B1 => n1880, B2 => n1611, C1 => n1437, C2 => 
                           n1950, A => n1004, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_18_port);
   U1450 : BUF_X1 port map( A => n976, Z => n1952);
   U1451 : BUF_X1 port map( A => n1876, Z => n1953);
   U1452 : NOR3_X1 port map( A1 => n1994, A2 => n109, A3 => n2095, ZN => n191);
   U1453 : BUF_X1 port map( A => n1863, Z => n1944);
   U1454 : INV_X1 port map( A => n1923, ZN => n1717);
   U1455 : AOI211_X1 port map( C1 => n1764, C2 => n1210, A => n882, B => n1641,
                           ZN => n916);
   U1456 : AOI211_X1 port map( C1 => n1635, C2 => n2076, A => n896, B => n1348,
                           ZN => n922);
   U1457 : NAND3_X1 port map( A1 => n1825, A2 => n1826, A3 => n1061, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_13_port);
   U1458 : AOI22_X1 port map( A1 => RF_WR_DATAx13x, A2 => n1948, B1 => 
                           RF_RD1_DATA(13), B2 => n1891, ZN => n1061);
   U1459 : OAI221_X1 port map( B1 => n1861, B2 => n1609, C1 => n1424, C2 => 
                           n1823, A => n1074, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_5_port);
   U1460 : INV_X1 port map( A => n1710, ZN => n441);
   U1461 : BUF_X2 port map( A => DATAPATH_IxThird_stxALU_IN2_1_port, Z => n1989
                           );
   U1462 : AND2_X1 port map( A1 => n887, A2 => n2073, ZN => n870);
   U1463 : AOI211_X1 port map( C1 => n1634, C2 => n2076, A => n896, B => n1347,
                           ZN => n921);
   U1464 : AOI211_X2 port map( C1 => n1706, C2 => n1298, A => n1995, B => n296,
                           ZN => n109);
   U1465 : INV_X1 port map( A => n785, ZN => n2145);
   U1466 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_1_port, ZN => 
                           n1574);
   U1467 : INV_X1 port map( A => n1574, ZN => n1575);
   U1468 : CLKBUF_X1 port map( A => n848, Z => n1576);
   U1469 : CLKBUF_X1 port map( A => n1942, Z => n1577);
   U1470 : CLKBUF_X3 port map( A => n1942, Z => n1578);
   U1471 : INV_X1 port map( A => n1862, ZN => n1942);
   U1472 : OR2_X1 port map( A1 => n1579, A2 => n1691, ZN => n831);
   U1473 : NOR2_X1 port map( A1 => n1712, A2 => n1916, ZN => n1579);
   U1474 : CLKBUF_X1 port map( A => n655, Z => n1580);
   U1475 : INV_X1 port map( A => n1651, ZN => n385);
   U1476 : XOR2_X1 port map( A => n1982, B => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, Z => n1651);
   U1477 : CLKBUF_X1 port map( A => n970, Z => n1581);
   U1478 : CLKBUF_X1 port map( A => n787, Z => n1582);
   U1479 : CLKBUF_X1 port map( A => n422, Z => n1583);
   U1480 : INV_X1 port map( A => n2137, ZN => n1584);
   U1481 : XNOR2_X1 port map( A => n2145, B => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, ZN => n1585);
   U1482 : CLKBUF_X1 port map( A => n742, Z => n1586);
   U1483 : INV_X2 port map( A => n1862, ZN => n1943);
   U1484 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_23_port, Z => 
                           n1587);
   U1485 : CLKBUF_X1 port map( A => n835, Z => n1875);
   U1486 : CLKBUF_X1 port map( A => n560, Z => n1588);
   U1487 : XNOR2_X1 port map( A => n1151, B => n1152, ZN => n1589);
   U1488 : BUF_X1 port map( A => n1689, Z => n1916);
   U1489 : INV_X1 port map( A => n108, ZN => n1819);
   U1490 : XNOR2_X1 port map( A => n1150, B => n1154, ZN => n1602);
   U1491 : OR2_X1 port map( A1 => n1865, A2 => n1335, ZN => n1603);
   U1492 : INV_X1 port map( A => n1729, ZN => n268);
   U1493 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_2_port, Z => n1988
                           );
   U1494 : AND3_X1 port map( A1 => n1128, A2 => n1127, A3 => n1126, ZN => n1623
                           );
   U1495 : AND3_X1 port map( A1 => n1104, A2 => n1103, A3 => n1102, ZN => n1624
                           );
   U1496 : AND3_X1 port map( A1 => n2112, A2 => n755, A3 => n597, ZN => n1631);
   U1497 : OR2_X1 port map( A1 => n1334, A2 => n1333, ZN => n1632);
   U1498 : INV_X1 port map( A => n1692, ZN => n647);
   U1499 : XNOR2_X1 port map( A => n1148, B => n1155, ZN => n1633);
   U1500 : BUF_X1 port map( A => n1601, Z => n1930);
   U1501 : AND3_X1 port map( A1 => n837, A2 => n152, A3 => n836, ZN => n1643);
   U1502 : AND3_X1 port map( A1 => n853, A2 => n180, A3 => n852, ZN => n1644);
   U1503 : CLKBUF_X1 port map( A => n953, Z => n1647);
   U1504 : AOI22_X1 port map( A1 => RF_WR_DATAx0x, A2 => n1948, B1 => 
                           RF_RD1_DATA(0), B2 => n1947, ZN => n1648);
   U1505 : INV_X1 port map( A => n1652, ZN => n446);
   U1506 : BUF_X1 port map( A => n985, Z => n1941);
   U1507 : AND2_X1 port map( A1 => n569, A2 => n1716, ZN => n1652);
   U1508 : AOI21_X1 port map( B1 => n1647, B2 => n808, A => n805, ZN => n1649);
   U1509 : CLKBUF_X1 port map( A => n518, Z => n1650);
   U1510 : INV_X2 port map( A => n1879, ZN => n1949);
   U1511 : NOR4_X1 port map( A1 => n1035, A2 => n1036, A3 => n333, A4 => n347, 
                           ZN => n1653);
   U1512 : NOR4_X1 port map( A1 => n1035, A2 => n1036, A3 => n333, A4 => n347, 
                           ZN => n1654);
   U1513 : NOR4_X1 port map( A1 => n1035, A2 => n1036, A3 => n333, A4 => n347, 
                           ZN => n969);
   U1514 : INV_X1 port map( A => n2113, ZN => n1655);
   U1515 : NAND2_X1 port map( A1 => n1732, A2 => n1733, ZN => n1656);
   U1516 : INV_X1 port map( A => n452, ZN => n1657);
   U1517 : XNOR2_X1 port map( A => n1658, B => n1929, ZN => n696);
   U1518 : XNOR2_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_0_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_0_port, ZN => n1658);
   U1519 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_3_port, Z => n1986
                           );
   U1520 : CLKBUF_X2 port map( A => DATAPATH_IxThird_stxALU_IN2_3_port, Z => 
                           n1987);
   U1521 : AND4_X1 port map( A1 => n1659, A2 => n1660, A3 => n1661, A4 => n1662
                           , ZN => n1094);
   U1522 : XNOR2_X1 port map( A => DATAPATH_IxWR_ADD_MEM_fu_4_port, B => n1893,
                           ZN => n1659);
   U1523 : XNOR2_X1 port map( A => n1147, B => n1163, ZN => n1660);
   U1524 : XOR2_X1 port map( A => DATAPATH_IxWR_ADD_MEM_fu_1_port, B => n1877, 
                           Z => n1661);
   U1525 : XOR2_X1 port map( A => n1813, B => n1151, Z => n1662);
   U1526 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_19_port, Z => 
                           n1663);
   U1527 : NAND2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN2_1_port, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, ZN => n1666);
   U1528 : NAND2_X1 port map( A1 => n1664, A2 => n1665, ZN => n1667);
   U1529 : NAND2_X1 port map( A1 => n1666, A2 => n1667, ZN => n1718);
   U1530 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_1_port, ZN => 
                           n1664);
   U1531 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_1_port, ZN => 
                           n1665);
   U1532 : OAI221_X1 port map( B1 => n1860, B2 => n1604, C1 => n1436, C2 => 
                           n1950, A => n1007, ZN => n1668);
   U1533 : OAI221_X1 port map( B1 => n1860, B2 => n1604, C1 => n1436, C2 => 
                           n1950, A => n1007, ZN => n1669);
   U1534 : INV_X1 port map( A => n2107, ZN => n1670);
   U1535 : OAI221_X1 port map( B1 => n1861, B2 => n1614, C1 => n1441, C2 => 
                           n1950, A => n988, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_22_port);
   U1536 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_21_port, Z => 
                           n1671);
   U1537 : CLKBUF_X1 port map( A => n594, Z => n1672);
   U1538 : XOR2_X1 port map( A => n2132, B => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, Z => n1673);
   U1539 : OAI221_X2 port map( B1 => n1860, B2 => n1607, C1 => n1448, C2 => 
                           n1951, A => n1032, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_29_port);
   U1540 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_25_port, Z => 
                           n1674);
   U1541 : OAI221_X1 port map( B1 => n1880, B2 => n1613, C1 => n1444, C2 => 
                           n1950, A => n1016, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_25_port);
   U1542 : AND4_X1 port map( A1 => n1653, A2 => n970, A3 => n968, A4 => n967, 
                           ZN => n1675);
   U1543 : AND4_X1 port map( A1 => n969, A2 => n970, A3 => n968, A4 => n967, ZN
                           => n1705);
   U1544 : NAND3_X1 port map( A1 => n1069, A2 => n1845, A3 => n1844, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_0_port);
   U1545 : OAI211_X1 port map( C1 => n1675, C2 => n1298, A => n1706, B => n1781
                           , ZN => n1676);
   U1546 : CLKBUF_X1 port map( A => n284, Z => n1677);
   U1547 : BUF_X1 port map( A => n1763, Z => n1764);
   U1548 : INV_X1 port map( A => n1158, ZN => RF_WR_ADD(4));
   U1549 : CLKBUF_X1 port map( A => n576, Z => n1679);
   U1550 : INV_X1 port map( A => n709, ZN => n1818);
   U1551 : INV_X1 port map( A => n713, ZN => n1817);
   U1552 : INV_X1 port map( A => n836, ZN => n1758);
   U1553 : INV_X1 port map( A => n1988, ZN => n1680);
   U1554 : INV_X2 port map( A => n1680, ZN => n1681);
   U1555 : NOR2_X1 port map( A1 => n2093, A2 => n1381, ZN => n1682);
   U1556 : NOR2_X1 port map( A1 => n2093, A2 => n1382, ZN => n1683);
   U1557 : NOR2_X1 port map( A1 => n2093, A2 => n1383, ZN => n1684);
   U1558 : NOR2_X1 port map( A1 => n2093, A2 => n1384, ZN => n1685);
   U1559 : NOR2_X1 port map( A1 => n2093, A2 => n1646, ZN => n1686);
   U1560 : NOR2_X1 port map( A1 => n2093, A2 => n1385, ZN => n1687);
   U1561 : NOR2_X1 port map( A1 => n1386, A2 => n2093, ZN => n1688);
   U1562 : AOI21_X1 port map( B1 => n819, B2 => n1689, A => n1690, ZN => n1691)
                           ;
   U1563 : OAI211_X1 port map( C1 => n1386, C2 => n1361, A => n833, B => n834, 
                           ZN => n819);
   U1564 : AND2_X1 port map( A1 => n658, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, ZN => n1692);
   U1565 : AND4_X1 port map( A1 => n1116, A2 => n1115, A3 => n1115, A4 => n1693
                           , ZN => n1808);
   U1566 : AOI22_X1 port map( A1 => RF_RD2_DATA(0), A2 => n985, B1 => n1577, B2
                           => RF_WR_DATAx0x, ZN => n1069);
   U1567 : AND4_X1 port map( A1 => n1633, A2 => n1602, A3 => n1694, A4 => n1589
                           , ZN => n1118);
   U1568 : INV_X1 port map( A => n1124, ZN => n1694);
   U1569 : AOI22_X1 port map( A1 => RF_RD2_DATA(3), A2 => n1808, B1 => n1578, 
                           B2 => RF_WR_DATAx3x, ZN => n1084);
   U1570 : NAND3_X1 port map( A1 => n1695, A2 => n1696, A3 => n1697, ZN => 
                           n1036);
   U1571 : INV_X1 port map( A => n642, ZN => n1695);
   U1572 : INV_X1 port map( A => n663, ZN => n1696);
   U1573 : INV_X1 port map( A => n624, ZN => n1697);
   U1574 : AND3_X1 port map( A1 => n1746, A2 => n1745, A3 => n1044, ZN => n2150
                           );
   U1575 : AND4_X2 port map( A1 => n1698, A2 => n1651, A3 => n1699, A4 => n1700
                           , ZN => n968);
   U1576 : INV_X1 port map( A => n371, ZN => n1698);
   U1577 : INV_X1 port map( A => n393, ZN => n1699);
   U1578 : INV_X1 port map( A => n1709, ZN => n1700);
   U1579 : NAND4_X1 port map( A1 => n1701, A2 => n1702, A3 => n1703, A4 => 
                           n1704, ZN => n1035);
   U1580 : INV_X1 port map( A => n686, ZN => n1701);
   U1581 : INV_X1 port map( A => n655, ZN => n1702);
   U1582 : INV_X1 port map( A => n353, ZN => n1703);
   U1583 : INV_X1 port map( A => n669, ZN => n1704);
   U1584 : OAI211_X1 port map( C1 => n1705, C2 => n1298, A => n1706, B => n1781
                           , ZN => n1780);
   U1585 : OAI21_X1 port map( B1 => n873, B2 => n874, A => n2072, ZN => n871);
   U1586 : INV_X1 port map( A => n899, ZN => n2072);
   U1587 : OAI22_X1 port map( A1 => n868, A2 => n869, B1 => n1353, B2 => n867, 
                           ZN => n181);
   U1588 : AND2_X1 port map( A1 => n1088, A2 => n2201, ZN => n979);
   U1589 : OAI211_X1 port map( C1 => n1386, C2 => n1361, A => n833, B => n834, 
                           ZN => n1712);
   U1590 : AND2_X1 port map( A1 => n1088, A2 => n2201, ZN => n1891);
   U1591 : AOI211_X1 port map( C1 => n706, C2 => n2101, A => n1335, B => n1337,
                           ZN => n703);
   U1592 : OAI22_X1 port map( A1 => n903, A2 => n904, B1 => n1707, B2 => n2070,
                           ZN => n876);
   U1593 : INV_X1 port map( A => n2057, ZN => n1708);
   U1594 : XOR2_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_0_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_0_port, Z => n1709);
   U1595 : XNOR2_X1 port map( A => n1921, B => n438, ZN => n1710);
   U1596 : INV_X1 port map( A => n1712, ZN => n1711);
   U1597 : CLKBUF_X1 port map( A => n469, Z => n1713);
   U1598 : OR2_X1 port map( A1 => n1870, A2 => n1628, ZN => n1714);
   U1599 : OR2_X1 port map( A1 => n1446, A2 => n1951, ZN => n1715);
   U1600 : NAND3_X1 port map( A1 => n1714, A2 => n1715, A3 => n1026, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_27_port);
   U1601 : BUF_X2 port map( A => n976, Z => n1951);
   U1602 : NAND3_X1 port map( A1 => n1648, A2 => n1728, A3 => n1727, ZN => 
                           n1716);
   U1603 : XNOR2_X1 port map( A => n1718, B => n1717, ZN => n568);
   U1604 : OR2_X1 port map( A1 => n1441, A2 => n1761, ZN => n1719);
   U1605 : OR2_X1 port map( A1 => n1179, A2 => n1769, ZN => n1720);
   U1606 : NAND3_X1 port map( A1 => n1719, A2 => n1720, A3 => n989, ZN => n747)
                           ;
   U1607 : CLKBUF_X1 port map( A => n618, Z => n1721);
   U1608 : OR2_X1 port map( A1 => n1435, A2 => n1762, ZN => n1722);
   U1609 : OR2_X1 port map( A1 => n1180, A2 => n1770, ZN => n1723);
   U1610 : NAND3_X1 port map( A1 => n1722, A2 => n1723, A3 => n992, ZN => n788)
                           ;
   U1611 : CLKBUF_X1 port map( A => n774, Z => n1724);
   U1612 : BUF_X2 port map( A => n1944, Z => n1769);
   U1613 : CLKBUF_X1 port map( A => n669, Z => n1725);
   U1614 : INV_X1 port map( A => n1764, ZN => n1726);
   U1615 : OR2_X1 port map( A1 => n1871, A2 => n1625, ZN => n1727);
   U1616 : OR2_X1 port map( A1 => n1419, A2 => n1823, ZN => n1728);
   U1617 : NAND3_X1 port map( A1 => n1068, A2 => n1728, A3 => n1727, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_0_port);
   U1618 : BUF_X2 port map( A => n1953, Z => n1871);
   U1619 : BUF_X2 port map( A => n1952, Z => n1823);
   U1620 : CLKBUF_X1 port map( A => n1755, Z => n1729);
   U1621 : OR2_X1 port map( A1 => n959, A2 => n1757, ZN => n1755);
   U1622 : NAND2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN2_2_port, A2 => 
                           n1731, ZN => n1732);
   U1623 : NAND2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_2_port, A2 => 
                           n1730, ZN => n1733);
   U1624 : NAND2_X1 port map( A1 => n1732, A2 => n1733, ZN => n438);
   U1625 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_2_port, ZN => 
                           n1730);
   U1626 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_2_port, ZN => 
                           n1731);
   U1627 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_2_port, Z => n1734
                           );
   U1628 : XNOR2_X1 port map( A => n2136, B => 
                           DATAPATH_IxThird_stxALU_IN1_26_port, ZN => n487);
   U1629 : CLKBUF_X1 port map( A => n2091, Z => n1735);
   U1630 : CLKBUF_X1 port map( A => n2134, Z => n1736);
   U1631 : OR2_X1 port map( A1 => n1447, A2 => n1761, ZN => n1737);
   U1632 : OR2_X1 port map( A1 => n1166, A2 => n1770, ZN => n1738);
   U1633 : NAND3_X1 port map( A1 => n1737, A2 => n1738, A3 => n1030, ZN => n735
                           );
   U1634 : XNOR2_X1 port map( A => n1986, B => n2126, ZN => n1739);
   U1635 : XNOR2_X1 port map( A => n1987, B => n2126, ZN => n1740);
   U1636 : OR2_X1 port map( A1 => n1422, A2 => n1761, ZN => n1741);
   U1637 : OR2_X1 port map( A1 => n1196, A2 => n1770, ZN => n1742);
   U1638 : NAND3_X1 port map( A1 => n1741, A2 => n1742, A3 => n1084, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_3_port);
   U1639 : BUF_X2 port map( A => n1944, Z => n1770);
   U1640 : CLKBUF_X1 port map( A => n568, Z => n1743);
   U1641 : CLKBUF_X2 port map( A => DATAPATH_IxThird_stxALU_IN2_0_port, Z => 
                           n1990);
   U1642 : OAI221_X4 port map( B1 => n1861, B2 => n1608, C1 => n1447, C2 => 
                           n1951, A => n1029, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_28_port);
   U1643 : CLKBUF_X1 port map( A => n779, Z => n1744);
   U1644 : OR2_X1 port map( A1 => n1433, A2 => n1762, ZN => n1745);
   U1645 : OR2_X1 port map( A1 => n1183, A2 => n1868, ZN => n1746);
   U1646 : NAND3_X1 port map( A1 => n1745, A2 => n1746, A3 => n1044, ZN => n760
                           );
   U1647 : OAI22_X1 port map( A1 => n2126, A2 => n778, B1 => n1744, B2 => n404,
                           ZN => n1747);
   U1648 : CLKBUF_X1 port map( A => n279, Z => n1748);
   U1649 : CLKBUF_X1 port map( A => n2102, Z => n1749);
   U1650 : CLKBUF_X1 port map( A => n1676, Z => n1750);
   U1651 : NAND2_X1 port map( A1 => n580, A2 => n1631, ZN => n754);
   U1652 : OAI22_X1 port map( A1 => n2122, A2 => n773, B1 => n1724, B2 => n359,
                           ZN => n1751);
   U1653 : NAND2_X1 port map( A1 => n181, A2 => n1644, ZN => n850);
   U1654 : NOR3_X1 port map( A1 => n1120, A2 => n1121, A3 => n1632, ZN => n1119
                           );
   U1655 : OR2_X1 port map( A1 => n1448, A2 => n1762, ZN => n1752);
   U1656 : OR2_X1 port map( A1 => n1157, A2 => n1868, ZN => n1753);
   U1657 : NAND3_X1 port map( A1 => n1752, A2 => n1753, A3 => n1033, ZN => n734
                           );
   U1658 : AND2_X1 port map( A1 => n1129, A2 => n1623, ZN => n1754);
   U1659 : NOR4_X2 port map( A1 => n1120, A2 => n1131, A3 => n1130, A4 => n1299
                           , ZN => n1129);
   U1660 : OR2_X1 port map( A1 => n1111, A2 => n1113, ZN => n1863);
   U1661 : OR2_X1 port map( A1 => n1875, A2 => n1916, ZN => n1756);
   U1662 : NAND2_X1 port map( A1 => n1756, A2 => n849, ZN => n848);
   U1663 : AND2_X1 port map( A1 => n1782, A2 => n1828, ZN => n1757);
   U1664 : XNOR2_X1 port map( A => n848, B => n1758, ZN => n1773);
   U1665 : CLKBUF_X1 port map( A => n282, Z => n1759);
   U1666 : CLKBUF_X1 port map( A => n1712, Z => n1760);
   U1667 : BUF_X2 port map( A => n981, Z => n1761);
   U1668 : BUF_X2 port map( A => n981, Z => n1762);
   U1669 : CLKBUF_X1 port map( A => n981, Z => n1945);
   U1670 : INV_X1 port map( A => n897, ZN => n1763);
   U1671 : AND2_X1 port map( A1 => n1676, A2 => CU_Ixcw2_i_12_port, ZN => n1772
                           );
   U1672 : CLKBUF_X1 port map( A => n897, Z => n1771);
   U1673 : INV_X1 port map( A => n1735, ZN => n1765);
   U1674 : CLKBUF_X1 port map( A => n766, Z => n1766);
   U1675 : CLKBUF_X1 port map( A => n758, Z => n1767);
   U1676 : CLKBUF_X1 port map( A => n696, Z => n1768);
   U1677 : AOI22_X1 port map( A1 => n897, A2 => n1368, B1 => n1772, B2 => n1378
                           , ZN => n283);
   U1678 : INV_X1 port map( A => n664, ZN => n1815);
   U1679 : NAND2_X1 port map( A1 => n835, A2 => n1643, ZN => n833);
   U1680 : CLKBUF_X1 port map( A => n815, Z => n1774);
   U1681 : CLKBUF_X1 port map( A => n1748, Z => n1775);
   U1682 : INV_X1 port map( A => n1750, ZN => n291);
   U1683 : CLKBUF_X1 port map( A => n745, Z => n1776);
   U1684 : CLKBUF_X1 port map( A => n738, Z => n1777);
   U1685 : OAI22_X1 port map( A1 => n1835, A2 => n765, B1 => n1766, B2 => n674,
                           ZN => n1778);
   U1686 : OAI22_X1 port map( A1 => n1979, A2 => n715, B1 => n716, B2 => n717, 
                           ZN => n1779);
   U1687 : OAI22_X1 port map( A1 => n1835, A2 => n765, B1 => n766, B2 => n674, 
                           ZN => n626);
   U1688 : XNOR2_X1 port map( A => n958, B => n1782, ZN => n815);
   U1689 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_30_port, Z => 
                           n1783);
   U1690 : INV_X1 port map( A => n2106, ZN => n1784);
   U1691 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_24_port, Z => 
                           n1785);
   U1692 : CLKBUF_X1 port map( A => n1716, Z => n1786);
   U1693 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_14_port, Z => 
                           n1787);
   U1694 : INV_X1 port map( A => n2049, ZN => n1788);
   U1695 : OR2_X1 port map( A1 => n1450, A2 => n1761, ZN => n1789);
   U1696 : OR2_X1 port map( A1 => n1170, A2 => n1769, ZN => n1790);
   U1697 : NAND3_X1 port map( A1 => n1789, A2 => n1790, A3 => n1014, ZN => n715
                           );
   U1698 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_4_port, Z => n1791
                           );
   U1699 : OR2_X1 port map( A1 => n1870, A2 => n1626, ZN => n1792);
   U1700 : OR2_X1 port map( A1 => n1430, A2 => n1951, ZN => n1793);
   U1701 : NAND3_X1 port map( A1 => n1792, A2 => n1793, A3 => n1057, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_11_port);
   U1702 : BUF_X1 port map( A => n1953, Z => n1870);
   U1703 : OAI221_X1 port map( B1 => n1861, B2 => n1606, C1 => n1428, C2 => 
                           n1951, A => n1040, ZN => n1794);
   U1704 : INV_X1 port map( A => n1001, ZN => n1795);
   U1705 : OAI221_X1 port map( B1 => n1861, B2 => n1597, C1 => n1435, C2 => 
                           n1950, A => n991, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_16_port);
   U1706 : BUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_12_port, Z => 
                           n1796);
   U1707 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_15_port, Z => 
                           n1797);
   U1708 : AND3_X2 port map( A1 => n1862, A2 => n1863, A3 => n1866, ZN => n985)
                           ;
   U1709 : CLKBUF_X1 port map( A => n551, Z => n1798);
   U1710 : OR2_X1 port map( A1 => n1440, A2 => n1761, ZN => n1799);
   U1711 : OR2_X1 port map( A1 => n1173, A2 => n1868, ZN => n1800);
   U1712 : NAND3_X1 port map( A1 => n1799, A2 => n1800, A3 => n998, ZN => n749)
                           ;
   U1713 : CLKBUF_X1 port map( A => n686, Z => n1801);
   U1714 : CLKBUF_X1 port map( A => n427, Z => n1802);
   U1715 : OR2_X1 port map( A1 => n1449, A2 => n1761, ZN => n1803);
   U1716 : OR2_X1 port map( A1 => n1169, A2 => n1869, ZN => n1804);
   U1717 : NAND3_X1 port map( A1 => n1803, A2 => n1804, A3 => n1011, ZN => n731
                           );
   U1718 : CLKBUF_X1 port map( A => n487, Z => n1805);
   U1719 : OR2_X1 port map( A1 => n1870, A2 => n1627, ZN => n1806);
   U1720 : OR2_X1 port map( A1 => n1445, A2 => n1951, ZN => n1807);
   U1721 : NAND3_X1 port map( A1 => n1806, A2 => n1807, A3 => n1023, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_26_port);
   U1722 : CLKBUF_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_8_port, Z => 
                           n1809);
   U1723 : OAI221_X1 port map( B1 => n1860, B2 => n1594, C1 => n1427, C2 => 
                           n1951, A => n1037, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_8_port);
   U1724 : XNOR2_X1 port map( A => n2365, B => n1164, ZN => n1107);
   U1725 : AND2_X1 port map( A1 => n1105, A2 => n1624, ZN => n1810);
   U1726 : INV_X1 port map( A => n1811, ZN => n1812);
   U1727 : XNOR2_X1 port map( A => DATAPATH_IxWR_ADD_MEM_fu_3_port, B => n1165,
                           ZN => n1097);
   U1728 : BUF_X1 port map( A => n976, Z => n1950);
   U1729 : AOI21_X1 port map( B1 => n1815, B2 => n626, A => n1692, ZN => n1814)
                           ;
   U1730 : BUF_X2 port map( A => n1808, Z => n1816);
   U1731 : XNOR2_X1 port map( A => DATAPATH_IxWR_ADD_MEM_fu_3_port, B => n1156,
                           ZN => n1121);
   U1732 : XNOR2_X1 port map( A => n1779, B => n1817, ZN => n712);
   U1733 : XNOR2_X1 port map( A => n708, B => n1818, ZN => n707);
   U1734 : OAI221_X1 port map( B1 => n1430, B2 => n1762, C1 => n1187, C2 => 
                           n1770, A => n1059, ZN => n1058);
   U1735 : OR4_X1 port map( A1 => n1994, A2 => n109, A3 => n159, A4 => n2094, 
                           ZN => n108);
   U1736 : AOI22_X1 port map( A1 => n1726, A2 => n1367, B1 => n1764, B2 => 
                           n1377, ZN => n1820);
   U1737 : OR2_X1 port map( A1 => n1429, A2 => n1945, ZN => n1821);
   U1738 : OR2_X1 port map( A1 => n1186, A2 => n1863, ZN => n1822);
   U1739 : NAND3_X1 port map( A1 => n1821, A2 => n1822, A3 => n1055, ZN => n768
                           );
   U1740 : CLKBUF_X1 port map( A => n294, Z => n1824);
   U1741 : OR2_X1 port map( A1 => n1861, A2 => n1630, ZN => n1825);
   U1742 : OR2_X1 port map( A1 => n1432, A2 => n1951, ZN => n1826);
   U1743 : CLKBUF_X1 port map( A => n903, Z => n1827);
   U1744 : AOI22_X1 port map( A1 => n1771, A2 => n1369, B1 => n1764, B2 => 
                           n1379, ZN => n1828);
   U1745 : AOI21_X1 port map( B1 => n1591, B2 => n2091, A => n279, ZN => n1829)
                           ;
   U1746 : OR2_X1 port map( A1 => n751, A2 => n582, ZN => n1830);
   U1747 : OR2_X1 port map( A1 => n2110, A2 => n753, ZN => n1831);
   U1748 : NAND3_X1 port map( A1 => n754, A2 => n1831, A3 => n1830, ZN => n520)
                           ;
   U1749 : OR2_X1 port map( A1 => n1860, A2 => n1629, ZN => n1832);
   U1750 : OR2_X1 port map( A1 => n1429, A2 => n1951, ZN => n1833);
   U1751 : NAND3_X1 port map( A1 => n1054, A2 => n1833, A3 => n1832, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_10_port);
   U1752 : NAND2_X1 port map( A1 => n1058, A2 => n1835, ZN => n1836);
   U1753 : NAND2_X1 port map( A1 => n1834, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, ZN => n1837);
   U1754 : NAND2_X1 port map( A1 => n1836, A2 => n1837, ZN => n669);
   U1755 : INV_X1 port map( A => n1058, ZN => n1834);
   U1756 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_11_port, ZN => 
                           n1835);
   U1757 : OAI22_X1 port map( A1 => n2115, A2 => n757, B1 => n1767, B2 => n630,
                           ZN => n1838);
   U1758 : OAI22_X1 port map( A1 => n2115, A2 => n757, B1 => n758, B2 => n630, 
                           ZN => n580);
   U1759 : OAI22_X1 port map( A1 => n1749, A2 => n737, B1 => n1777, B2 => n475,
                           ZN => n1839);
   U1760 : CLKBUF_X1 port map( A => n1747, Z => n1840);
   U1761 : OAI22_X1 port map( A1 => n2126, A2 => n778, B1 => n779, B2 => n404, 
                           ZN => n357);
   U1762 : INV_X1 port map( A => n1892, ZN => n1841);
   U1763 : INV_X1 port map( A => n1849, ZN => n1842);
   U1764 : XOR2_X1 port map( A => n1736, B => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, Z => n1843);
   U1765 : OR2_X1 port map( A1 => n1419, A2 => n1945, ZN => n1844);
   U1766 : OR2_X1 port map( A1 => n1193, A2 => n1863, ZN => n1845);
   U1767 : BUF_X2 port map( A => n1944, Z => n1868);
   U1768 : OAI22_X1 port map( A1 => n2106, A2 => n744, B1 => n1776, B2 => n524,
                           ZN => n1846);
   U1769 : OAI22_X1 port map( A1 => n2106, A2 => n744, B1 => n745, B2 => n524, 
                           ZN => n471);
   U1770 : CLKBUF_X1 port map( A => n353, Z => n1847);
   U1771 : OAI22_X1 port map( A1 => n1383, A2 => n1636, B1 => n1649, B2 => n799
                           , ZN => n1848);
   U1772 : OAI22_X1 port map( A1 => n1383, A2 => n1636, B1 => n952, B2 => n799,
                           ZN => n936);
   U1773 : CLKBUF_X1 port map( A => n326, Z => n1849);
   U1774 : CLKBUF_X1 port map( A => n868, Z => n1850);
   U1775 : OAI22_X1 port map( A1 => n1346, A2 => n2079, B1 => n929, B2 => n930,
                           ZN => n919);
   U1776 : NAND2_X1 port map( A1 => n1129, A2 => n1623, ZN => n1115);
   U1777 : CLKBUF_X1 port map( A => n1839, Z => n1851);
   U1778 : OAI22_X1 port map( A1 => n1749, A2 => n737, B1 => n738, B2 => n475, 
                           ZN => n429);
   U1779 : CLKBUF_X1 port map( A => n520, Z => n1852);
   U1780 : NOR4_X1 port map( A1 => n560, A2 => n576, A3 => n536, A4 => n618, ZN
                           => n1856);
   U1781 : AND4_X1 port map( A1 => n1853, A2 => n1854, A3 => n1856, A4 => n1855
                           , ZN => n970);
   U1782 : AND4_X1 port map( A1 => n1022, A2 => BRANCH_EN_i, A3 => n463, A4 => 
                           n1673, ZN => n1853);
   U1783 : NOR4_X1 port map( A1 => n512, A2 => n503, A3 => n427, A4 => n422, ZN
                           => n1854);
   U1784 : NOR4_X1 port map( A1 => n610, A2 => n1585, A3 => n518, A4 => n551, 
                           ZN => n1855);
   U1785 : OAI22_X1 port map( A1 => n1707, A2 => n2070, B1 => n1827, B2 => n904
                           , ZN => n1857);
   U1786 : BUF_X2 port map( A => n1944, Z => n1869);
   U1787 : CLKBUF_X1 port map( A => n1930, Z => n1929);
   U1788 : CLKBUF_X1 port map( A => n1922, Z => n1928);
   U1789 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_5_port, ZN => 
                           n1982);
   U1790 : NAND2_X1 port map( A1 => n1105, A2 => n1624, ZN => n1093);
   U1791 : OAI22_X1 port map( A1 => n1353, A2 => n867, B1 => n1850, B2 => n869,
                           ZN => n1858);
   U1792 : OAI22_X1 port map( A1 => n1353, A2 => n867, B1 => n1850, B2 => n869,
                           ZN => n1859);
   U1793 : BUF_X2 port map( A => n1953, Z => n1860);
   U1794 : BUF_X2 port map( A => n1953, Z => n1861);
   U1795 : NOR2_X1 port map( A1 => n1912, A2 => n1921, ZN => n401);
   U1796 : INV_X1 port map( A => n571, ZN => n2160);
   U1797 : XNOR2_X1 port map( A => n709, B => n717, ZN => n726);
   U1798 : XNOR2_X1 port map( A => n713, B => n717, ZN => n725);
   U1799 : INV_X1 port map( A => n882, ZN => n2076);
   U1800 : INV_X1 port map( A => n1930, ZN => n1920);
   U1801 : INV_X1 port map( A => n1930, ZN => n1919);
   U1802 : INV_X1 port map( A => n1930, ZN => n1921);
   U1803 : BUF_X1 port map( A => n1978, Z => n1873);
   U1804 : BUF_X1 port map( A => n1978, Z => n1872);
   U1805 : INV_X1 port map( A => n1929, ZN => n1918);
   U1806 : AOI21_X1 port map( B1 => n405, B2 => n406, A => n407, ZN => n403);
   U1807 : XNOR2_X1 port map( A => n1918, B => n1657, ZN => n454);
   U1808 : BUF_X1 port map( A => n108, Z => n1903);
   U1809 : BUF_X1 port map( A => n299, Z => n1962);
   U1810 : BUF_X1 port map( A => n108, Z => n1901);
   U1811 : BUF_X1 port map( A => n2013, Z => n1905);
   U1812 : BUF_X1 port map( A => n108, Z => n1902);
   U1813 : BUF_X1 port map( A => n54, Z => n1966);
   U1814 : BUF_X1 port map( A => n54, Z => n1967);
   U1815 : BUF_X1 port map( A => n299, Z => n1961);
   U1816 : BUF_X1 port map( A => n2013, Z => n1904);
   U1817 : BUF_X1 port map( A => n2014, Z => n1907);
   U1818 : BUF_X1 port map( A => n2014, Z => n1906);
   U1819 : BUF_X1 port map( A => n54, Z => n1968);
   U1820 : AOI21_X1 port map( B1 => n364, B2 => n361, A => n362, ZN => n363);
   U1821 : AOI21_X1 port map( B1 => n360, B2 => n361, A => n362, ZN => n358);
   U1822 : AOI21_X1 port map( B1 => n587, B2 => n584, A => n585, ZN => n586);
   U1823 : INV_X1 port map( A => n783, ZN => n2112);
   U1824 : INV_X1 port map( A => n464, ZN => n2100);
   U1825 : BUF_X1 port map( A => n2162, Z => n1912);
   U1826 : BUF_X1 port map( A => n2162, Z => n1911);
   U1827 : AOI21_X1 port map( B1 => n412, B2 => n406, A => n407, ZN => n411);
   U1828 : AOI21_X1 port map( B1 => n635, B2 => n632, A => n633, ZN => n634);
   U1829 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n633, ZN => n629);
   U1830 : NOR2_X1 port map( A1 => n1929, A2 => n1912, ZN => n571);
   U1831 : XNOR2_X1 port map( A => n405, B => n441, ZN => n440);
   U1832 : BUF_X1 port map( A => n1978, Z => n1874);
   U1833 : BUF_X1 port map( A => n2162, Z => n1913);
   U1834 : INV_X1 port map( A => n1977, ZN => n1969);
   U1835 : INV_X1 port map( A => n1977, ZN => n1970);
   U1836 : INV_X1 port map( A => n1938, ZN => n1931);
   U1837 : XNOR2_X1 port map( A => n870, B => n886, ZN => n889);
   U1838 : XNOR2_X1 port map( A => n870, B => n885, ZN => n890);
   U1839 : XNOR2_X1 port map( A => n1924, B => n1788, ZN => n717);
   U1840 : OAI211_X1 port map( C1 => n2160, C2 => n562, A => n563, B => n564, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_1_port);
   U1841 : XNOR2_X1 port map( A => n446, B => n1743, ZN => n562);
   U1842 : AOI22_X1 port map( A1 => n2128, A2 => n1989, B1 => n401, B2 => n567,
                           ZN => n563);
   U1843 : NOR2_X1 port map( A1 => n365, A2 => n2123, ZN => n362);
   U1844 : NOR2_X1 port map( A1 => n588, A2 => n2111, ZN => n585);
   U1845 : XNOR2_X1 port map( A => n1927, B => n624, ZN => n630);
   U1846 : XNOR2_X1 port map( A => n1924, B => n1713, ZN => n475);
   U1847 : XNOR2_X1 port map( A => n1919, B => n371, ZN => n375);
   U1848 : XNOR2_X1 port map( A => n1986, B => n2126, ZN => n399);
   U1849 : AOI21_X1 port map( B1 => n432, B2 => n727, A => n719, ZN => n709);
   U1850 : AOI21_X1 port map( B1 => n434, B2 => n727, A => n719, ZN => n713);
   U1851 : XNOR2_X1 port map( A => n1922, B => n1986, ZN => n778);
   U1852 : OAI21_X1 port map( B1 => n568, B2 => n781, A => n444, ZN => n780);
   U1853 : OAI21_X1 port map( B1 => n776, B2 => n387, A => n378, ZN => n775);
   U1854 : INV_X1 port map( A => n379, ZN => n2124);
   U1855 : BUF_X1 port map( A => n92, Z => n1963);
   U1856 : BUF_X1 port map( A => n92, Z => n1964);
   U1857 : BUF_X1 port map( A => n2005, Z => n1899);
   U1858 : BUF_X1 port map( A => n2005, Z => n1898);
   U1859 : NOR2_X1 port map( A1 => n530, A2 => n2107, ZN => n527);
   U1860 : NOR2_X1 port map( A1 => n636, A2 => n2116, ZN => n633);
   U1861 : OAI21_X1 port map( B1 => n442, B2 => n443, A => n444, ZN => n405);
   U1862 : NOR2_X1 port map( A1 => n680, A2 => n2118, ZN => n677);
   U1863 : BUF_X1 port map( A => n2005, Z => n1900);
   U1864 : NOR2_X1 port map( A1 => n413, A2 => n2127, ZN => n407);
   U1865 : NOR2_X1 port map( A1 => n481, A2 => n2103, ZN => n478);
   U1866 : XNOR2_X1 port map( A => n1928, B => n1847, ZN => n359);
   U1867 : XNOR2_X1 port map( A => n1920, B => 
                           DATAPATH_IxThird_stxALU_IN2_1_port, ZN => n447);
   U1868 : XNOR2_X1 port map( A => n1920, B => n1980, ZN => n380);
   U1869 : OAI21_X1 port map( B1 => n1814, B2 => n657, A => n648, ZN => n759);
   U1870 : AOI22_X1 port map( A1 => n613, A2 => n2113, B1 => n2148, B2 => n2114
                           , ZN => n611);
   U1871 : XNOR2_X1 port map( A => n1925, B => n503, ZN => n505);
   U1872 : AOI22_X1 port map( A1 => n1908, A2 => n371, B1 => 
                           DATAPATH_IxThird_stxALU1xN197, B2 => n1960, ZN => 
                           n370);
   U1873 : XNOR2_X1 port map( A => n1923, B => n385, ZN => n387);
   U1874 : INV_X1 port map( A => n190, ZN => n2014);
   U1875 : OAI21_X1 port map( B1 => n377, B2 => n379, A => n378, ZN => n364);
   U1876 : OAI21_X1 port map( B1 => n376, B2 => n377, A => n378, ZN => n360);
   U1877 : XNOR2_X1 port map( A => n1919, B => n347, ZN => n348);
   U1878 : INV_X1 port map( A => n191, ZN => n2013);
   U1879 : XNOR2_X1 port map( A => n1918, B => n512, ZN => n513);
   U1880 : XNOR2_X1 port map( A => n1920, B => n393, ZN => n394);
   U1881 : NOR2_X1 port map( A1 => n582, A2 => n619, ZN => n755);
   U1882 : AOI21_X1 port map( B1 => n2125, B2 => n379, A => n376, ZN => n386);
   U1883 : NAND2_X1 port map( A1 => n1991, A2 => n1963, ZN => n299);
   U1884 : NAND2_X1 port map( A1 => n1900, A2 => n1991, ZN => n54);
   U1885 : INV_X1 port map( A => n601, ZN => n2148);
   U1886 : INV_X1 port map( A => CU_IxN25, ZN => n1999);
   U1887 : OAI211_X1 port map( C1 => n395, C2 => n2160, A => n397, B => n398, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_3_port);
   U1888 : XNOR2_X1 port map( A => n404, B => n411, ZN => n395);
   U1889 : AOI22_X1 port map( A1 => n400, A2 => n1987, B1 => n401, B2 => n402, 
                           ZN => n397);
   U1890 : AOI22_X1 port map( A1 => n1908, A2 => n1740, B1 => 
                           DATAPATH_IxThird_stxALU1xN194, B2 => n1960, ZN => 
                           n398);
   U1891 : INV_X1 port map( A => n729, ZN => n2133);
   U1892 : OAI211_X1 port map( C1 => n435, C2 => n2160, A => n436, B => n437, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_2_port);
   U1893 : XNOR2_X1 port map( A => n412, B => n1710, ZN => n435);
   U1894 : AOI22_X1 port map( A1 => n439, A2 => n1681, B1 => n401, B2 => n440, 
                           ZN => n436);
   U1895 : AOI22_X1 port map( A1 => n1908, A2 => n1656, B1 => 
                           DATAPATH_IxThird_stxALU1xN193, B2 => n1960, ZN => 
                           n437);
   U1896 : XNOR2_X1 port map( A => n1918, B => n2135, ZN => n737);
   U1897 : OAI21_X1 port map( B1 => n740, B2 => n505, A => n492, ZN => n739);
   U1898 : NOR2_X1 port map( A1 => n2203, A2 => n1902, ZN => n168);
   U1899 : NAND2_X1 port map( A1 => n2065, A2 => n2071, ZN => n900);
   U1900 : BUF_X1 port map( A => n1927, Z => n1924);
   U1901 : BUF_X1 port map( A => n92, Z => n1965);
   U1902 : NAND2_X1 port map( A1 => n600, A2 => n602, ZN => n587);
   U1903 : OR3_X1 port map( A1 => n599, A2 => n2113, A3 => n2148, ZN => n602);
   U1904 : INV_X1 port map( A => n103, ZN => n2012);
   U1905 : BUF_X1 port map( A => n1930, Z => n1922);
   U1906 : BUF_X1 port map( A => n1601, Z => n1923);
   U1907 : BUF_X1 port map( A => n1930, Z => n1927);
   U1908 : INV_X1 port map( A => n1997, ZN => CU_Ixcw_LUT_6_port);
   U1909 : INV_X1 port map( A => n732, ZN => n2098);
   U1910 : BUF_X1 port map( A => n1930, Z => n1926);
   U1911 : INV_X1 port map( A => n182, ZN => n2050);
   U1912 : INV_X1 port map( A => n46, ZN => n2054);
   U1913 : INV_X1 port map( A => n48, ZN => n2085);
   U1914 : INV_X1 port map( A => n49, ZN => n2090);
   U1915 : INV_X1 port map( A => n1979, ZN => n1978);
   U1916 : INV_X1 port map( A => n217, ZN => n2068);
   U1917 : INV_X1 port map( A => n206, ZN => n2066);
   U1918 : INV_X1 port map( A => n1603, ZN => n1954);
   U1919 : INV_X1 port map( A => n1603, ZN => n1955);
   U1920 : OAI21_X1 port map( B1 => n443, B2 => n446, A => n444, ZN => n412);
   U1921 : BUF_X1 port map( A => n2159, Z => n1908);
   U1922 : OAI21_X1 port map( B1 => n646, B2 => n647, A => n648, ZN => n631);
   U1923 : OAI21_X1 port map( B1 => n649, B2 => n646, A => n648, ZN => n635);
   U1924 : AOI21_X1 port map( B1 => n679, B2 => n676, A => n677, ZN => n678);
   U1925 : AOI21_X1 port map( B1 => n529, B2 => n526, A => n527, ZN => n528);
   U1926 : AOI21_X1 port map( B1 => n583, B2 => n584, A => n585, ZN => n581);
   U1927 : AOI21_X1 port map( B1 => n675, B2 => n676, A => n677, ZN => n673);
   U1928 : AOI21_X1 port map( B1 => n480, B2 => n477, A => n478, ZN => n479);
   U1929 : AOI21_X1 port map( B1 => n476, B2 => n477, A => n478, ZN => n474);
   U1930 : BUF_X1 port map( A => n2159, Z => n1909);
   U1931 : AOI21_X1 port map( B1 => n525, B2 => n526, A => n527, ZN => n523);
   U1932 : BUF_X1 port map( A => n2159, Z => n1910);
   U1933 : NAND2_X1 port map( A1 => n530, A2 => n2107, ZN => n526);
   U1934 : NAND2_X1 port map( A1 => n588, A2 => n2111, ZN => n584);
   U1935 : NAND2_X1 port map( A1 => n636, A2 => n2116, ZN => n632);
   U1936 : NAND2_X1 port map( A1 => n413, A2 => n2127, ZN => n406);
   U1937 : NAND2_X1 port map( A1 => n365, A2 => n2123, ZN => n361);
   U1938 : NAND2_X1 port map( A1 => n680, A2 => n2118, ZN => n676);
   U1939 : NAND2_X1 port map( A1 => n481, A2 => n2103, ZN => n477);
   U1940 : INV_X1 port map( A => n421, ZN => n2162);
   U1941 : INV_X1 port map( A => n28, ZN => n2004);
   U1942 : BUF_X1 port map( A => n1930, Z => n1925);
   U1943 : INV_X1 port map( A => n1797, ZN => n2115);
   U1944 : XNOR2_X1 port map( A => n1919, B => n2149, ZN => n757);
   U1945 : NAND2_X1 port map( A1 => n2073, A2 => n884, ZN => n879);
   U1946 : NOR2_X1 port map( A1 => n270, A2 => n271, ZN => n269);
   U1947 : INV_X1 port map( A => n109, ZN => n2015);
   U1948 : XNOR2_X1 port map( A => n861, B => n855, ZN => n857);
   U1949 : XNOR2_X1 port map( A => n851, B => n855, ZN => n858);
   U1950 : OAI21_X1 port map( B1 => n1917, B2 => n1639, A => n862, ZN => n861);
   U1951 : OAI21_X1 port map( B1 => n941, B2 => n946, A => n2195, ZN => n944);
   U1952 : XNOR2_X1 port map( A => n844, B => n839, ZN => n840);
   U1953 : XNOR2_X1 port map( A => n834, B => n839, ZN => n841);
   U1954 : OAI21_X1 port map( B1 => n1917, B2 => n1640, A => n845, ZN => n844);
   U1955 : OAI21_X1 port map( B1 => n804, B2 => n801, A => n2198, ZN => n803);
   U1956 : INV_X1 port map( A => n1982, ZN => n1980);
   U1957 : XNOR2_X1 port map( A => n1920, B => n771, ZN => n337);
   U1958 : XNOR2_X1 port map( A => n1920, B => n1586, ZN => n495);
   U1959 : OAI21_X1 port map( B1 => n1135, B2 => n2043, A => n1134, ZN => 
                           CU_IxN25);
   U1960 : INV_X1 port map( A => n27, ZN => n2043);
   U1961 : AOI21_X1 port map( B1 => n1137, B2 => n2045, A => n1138, ZN => n1135
                           );
   U1962 : XNOR2_X1 port map( A => n372, B => n2123, ZN => n371);
   U1963 : XNOR2_X1 port map( A => n1918, B => n735, ZN => n457);
   U1964 : NAND2_X1 port map( A1 => n877, A2 => n900, ZN => n898);
   U1965 : XNOR2_X1 port map( A => n1919, B => n1834, ZN => n765);
   U1966 : XNOR2_X1 port map( A => n789, B => n2102, ZN => n469);
   U1967 : XNOR2_X1 port map( A => n2155, B => 
                           DATAPATH_IxThird_stxALU_IN1_8_port, ZN => n347);
   U1968 : XNOR2_X1 port map( A => n2156, B => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, ZN => n353);
   U1969 : XNOR2_X1 port map( A => n1985, B => 
                           DATAPATH_IxThird_stxALU_IN1_4_port, ZN => n393);
   U1970 : AOI21_X1 port map( B1 => n101, B2 => n1819, A => n109, ZN => n103);
   U1971 : AOI21_X1 port map( B1 => n132, B2 => n1819, A => n109, ZN => n139);
   U1972 : AOI21_X1 port map( B1 => n144, B2 => n1819, A => n109, ZN => n150);
   U1973 : AOI21_X1 port map( B1 => n172, B2 => n1819, A => n109, ZN => n179);
   U1974 : AOI21_X1 port map( B1 => n198, B2 => n1819, A => n109, ZN => n205);
   U1975 : XNOR2_X1 port map( A => n1918, B => n734, ZN => n729);
   U1976 : XNOR2_X1 port map( A => n2149, B => 
                           DATAPATH_IxThird_stxALU_IN1_15_port, ZN => n624);
   U1977 : AOI21_X1 port map( B1 => n1957, B2 => n1670, A => n1955, ZN => n534)
                           ;
   U1978 : INV_X1 port map( A => n1583, ZN => n2049);
   U1979 : AOI21_X1 port map( B1 => n1957, B2 => n1872, A => n1954, ZN => n416)
                           ;
   U1980 : AOI22_X1 port map( A1 => n1872, A2 => n1958, B1 => n420, B2 => n421,
                           ZN => n419);
   U1981 : XNOR2_X1 port map( A => n1919, B => n2156, ZN => n773);
   U1982 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_7_port, ZN => 
                           n2122);
   U1983 : AOI21_X1 port map( B1 => n775, B2 => n375, A => n362, ZN => n774);
   U1984 : NAND2_X1 port map( A1 => n912, A2 => n2067, ZN => n927);
   U1985 : INV_X1 port map( A => n921, ZN => n2067);
   U1986 : OAI22_X1 port map( A1 => n2097, A2 => n2133, B1 => n722, B2 => n454,
                           ZN => n718);
   U1987 : OAI221_X1 port map( B1 => n1911, B2 => n590, C1 => n2145, C2 => n592
                           , A => n593, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_18_port);
   U1988 : AOI21_X1 port map( B1 => n1956, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, A => n1955, ZN 
                           => n592);
   U1989 : INV_X1 port map( A => n965, ZN => n2092);
   U1990 : AOI21_X1 port map( B1 => n962, B2 => n961, A => n1386, ZN => n965);
   U1991 : OAI221_X1 port map( B1 => n2137, B2 => n500, C1 => n1912, C2 => n501
                           , A => n502, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_25_port);
   U1992 : AOI21_X1 port map( B1 => n1957, B2 => n1674, A => n1955, ZN => n500)
                           ;
   U1993 : AOI22_X1 port map( A1 => n1909, A2 => n503, B1 => 
                           DATAPATH_IxThird_stxALU1xN216, B2 => n1959, ZN => 
                           n502);
   U1994 : XNOR2_X1 port map( A => n2154, B => 
                           DATAPATH_IxThird_stxALU_IN1_9_port, ZN => n333);
   U1995 : OAI221_X1 port map( B1 => n1911, B2 => n349, C1 => n2156, C2 => n351
                           , A => n352, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_7_port);
   U1996 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, A => n1954, ZN 
                           => n351);
   U1997 : AOI22_X1 port map( A1 => n1908, A2 => n1847, B1 => 
                           DATAPATH_IxThird_stxALU1xN198, B2 => n1960, ZN => 
                           n352);
   U1998 : OAI221_X1 port map( B1 => n1911, B2 => n367, C1 => n2157, C2 => n369
                           , A => n370, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_6_port);
   U1999 : INV_X1 port map( A => n372, ZN => n2157);
   U2000 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_6_port, A => n1954, ZN 
                           => n369);
   U2001 : OAI221_X1 port map( B1 => n1911, B2 => n423, C1 => n2131, C2 => n425
                           , A => n426, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_30_port);
   U2002 : AOI21_X1 port map( B1 => n1957, B2 => n1783, A => n1954, ZN => n425)
                           ;
   U2003 : OAI221_X1 port map( B1 => n1911, B2 => n620, C1 => n2149, C2 => n622
                           , A => n623, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_15_port);
   U2004 : AOI21_X1 port map( B1 => n1957, B2 => n1797, A => n1955, ZN => n622)
                           ;
   U2005 : AOI22_X1 port map( A1 => n1910, A2 => n624, B1 => 
                           DATAPATH_IxThird_stxALU1xN206, B2 => n1958, ZN => 
                           n623);
   U2006 : OAI221_X1 port map( B1 => n1911, B2 => n638, C1 => n2150, C2 => n640
                           , A => n641, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_14_port);
   U2007 : AOI21_X1 port map( B1 => n1956, B2 => n1787, A => n1954, ZN => n640)
                           ;
   U2008 : OAI221_X1 port map( B1 => n1736, B2 => n459, C1 => n1912, C2 => n460
                           , A => n461, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_28_port);
   U2009 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, A => n1954, ZN 
                           => n459);
   U2010 : AOI22_X1 port map( A1 => n1908, A2 => n2099, B1 => 
                           DATAPATH_IxThird_stxALU1xN219, B2 => n1959, ZN => 
                           n461);
   U2011 : XNOR2_X1 port map( A => n2101, B => n464, ZN => n460);
   U2012 : OAI221_X1 port map( B1 => n1911, B2 => n465, C1 => n2135, C2 => n467
                           , A => n468, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_27_port);
   U2013 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_27_port, A => n1954, ZN 
                           => n467);
   U2014 : AOI22_X1 port map( A1 => n1908, A2 => n1713, B1 => 
                           DATAPATH_IxThird_stxALU1xN218, B2 => n1959, ZN => 
                           n468);
   U2015 : OAI221_X1 port map( B1 => n1911, B2 => n483, C1 => n2136, C2 => n485
                           , A => n486, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_26_port);
   U2016 : INV_X1 port map( A => n488, ZN => n2136);
   U2017 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_26_port, A => n1954, ZN 
                           => n485);
   U2018 : AOI22_X1 port map( A1 => n1909, A2 => n1805, B1 => 
                           DATAPATH_IxThird_stxALU1xN217, B2 => n1959, ZN => 
                           n486);
   U2019 : OAI221_X1 port map( B1 => n2132, B2 => n449, C1 => n1912, C2 => n450
                           , A => n451, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_29_port);
   U2020 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, A => n1954, ZN 
                           => n449);
   U2021 : AOI22_X1 port map( A1 => n1908, A2 => n452, B1 => 
                           DATAPATH_IxThird_stxALU1xN220, B2 => n1959, ZN => 
                           n451);
   U2022 : XNOR2_X1 port map( A => n453, B => n454, ZN => n450);
   U2023 : OAI221_X1 port map( B1 => n2138, B2 => n509, C1 => n1912, C2 => n510
                           , A => n511, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_24_port);
   U2024 : AOI21_X1 port map( B1 => n1957, B2 => n1785, A => n1955, ZN => n509)
                           ;
   U2025 : AOI22_X1 port map( A1 => n1909, A2 => n512, B1 => 
                           DATAPATH_IxThird_stxALU1xN215, B2 => n1959, ZN => 
                           n511);
   U2026 : OAI221_X1 port map( B1 => n2152, B2 => n660, C1 => n1912, C2 => n661
                           , A => n662, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_12_port);
   U2027 : AOI21_X1 port map( B1 => n1956, B2 => n1796, A => n1954, ZN => n660)
                           ;
   U2028 : AOI22_X1 port map( A1 => n1910, A2 => n663, B1 => 
                           DATAPATH_IxThird_stxALU1xN203, B2 => n1958, ZN => 
                           n662);
   U2029 : OAI221_X1 port map( B1 => n1911, B2 => n665, C1 => n1834, C2 => n667
                           , A => n668, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_11_port);
   U2030 : AOI21_X1 port map( B1 => n1956, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, A => n1954, ZN 
                           => n667);
   U2031 : OAI221_X1 port map( B1 => n2154, B2 => n328, C1 => n1912, C2 => n330
                           , A => n331, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_9_port);
   U2032 : AOI21_X1 port map( B1 => n1956, B2 => n1794, A => n1954, ZN => n328)
                           ;
   U2033 : AOI22_X1 port map( A1 => n1908, A2 => n333, B1 => 
                           DATAPATH_IxThird_stxALU1xN200, B2 => n1958, ZN => 
                           n331);
   U2034 : XNOR2_X1 port map( A => n335, B => n336, ZN => n330);
   U2035 : OAI221_X1 port map( B1 => n2155, B2 => n344, C1 => n1913, C2 => n345
                           , A => n346, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_8_port);
   U2036 : AOI21_X1 port map( B1 => n1957, B2 => n1809, A => n1954, ZN => n344)
                           ;
   U2037 : AOI22_X1 port map( A1 => n1908, A2 => n347, B1 => 
                           DATAPATH_IxThird_stxALU1xN199, B2 => n1960, ZN => 
                           n346);
   U2038 : OAI221_X1 port map( B1 => n1912, B2 => n682, C1 => n2153, C2 => n684
                           , A => n685, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_10_port);
   U2039 : AOI21_X1 port map( B1 => n1956, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, A => n1954, ZN 
                           => n684);
   U2040 : OAI221_X1 port map( B1 => n2143, B2 => n557, C1 => n1912, C2 => n558
                           , A => n559, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_20_port);
   U2041 : AOI21_X1 port map( B1 => n1956, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, A => n1955, ZN 
                           => n557);
   U2042 : OAI221_X1 port map( B1 => n1985, B2 => n390, C1 => n1913, C2 => n391
                           , A => n392, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_4_port);
   U2043 : AOI21_X1 port map( B1 => n1957, B2 => n1791, A => n1954, ZN => n390)
                           ;
   U2044 : AOI22_X1 port map( A1 => n1908, A2 => n393, B1 => 
                           DATAPATH_IxThird_stxALU1xN195, B2 => n1960, ZN => 
                           n392);
   U2045 : INV_X1 port map( A => n340, ZN => n2120);
   U2046 : AOI21_X1 port map( B1 => n911, B2 => n921, A => n922, ZN => n910);
   U2047 : AND2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_28_port, A2 => 
                           n457, ZN => n455);
   U2048 : OAI221_X1 port map( B1 => n2151, B2 => n652, C1 => n1912, C2 => n653
                           , A => n654, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_13_port);
   U2049 : AOI21_X1 port map( B1 => n1956, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, A => n1954, ZN 
                           => n652);
   U2050 : AOI22_X1 port map( A1 => n1910, A2 => n1580, B1 => 
                           DATAPATH_IxThird_stxALU1xN204, B2 => n1958, ZN => 
                           n654);
   U2051 : XNOR2_X1 port map( A => n2152, B => 
                           DATAPATH_IxThird_stxALU_IN1_12_port, ZN => n663);
   U2052 : OAI221_X1 port map( B1 => n1982, B2 => n382, C1 => n1913, C2 => n383
                           , A => n384, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_5_port);
   U2053 : AOI21_X1 port map( B1 => n1957, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, A => n1954, ZN 
                           => n382);
   U2054 : AOI22_X1 port map( A1 => n1908, A2 => n385, B1 => 
                           DATAPATH_IxThird_stxALU1xN196, B2 => n1960, ZN => 
                           n384);
   U2055 : AOI21_X1 port map( B1 => n2109, B2 => n2144, A => n555, ZN => n552);
   U2056 : INV_X1 port map( A => n543, ZN => n2144);
   U2057 : INV_X1 port map( A => n1451, ZN => n2093);
   U2058 : XNOR2_X1 port map( A => n2132, B => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, ZN => n452);
   U2059 : XNOR2_X1 port map( A => n1924, B => n372, ZN => n365);
   U2060 : OR2_X2 port map( A1 => n2200, A2 => n1111, ZN => n1862);
   U2061 : NOR3_X1 port map( A1 => IRAM_ADD_23_port, A2 => n144, A3 => n1902, 
                           ZN => n156);
   U2062 : XNOR2_X1 port map( A => n1928, B => n768, ZN => n680);
   U2063 : XNOR2_X1 port map( A => n1918, B => n1584, ZN => n498);
   U2064 : XNOR2_X1 port map( A => n1925, B => n488, ZN => n481);
   U2065 : AOI21_X1 port map( B1 => n809, B2 => n2084, A => n811, ZN => n800);
   U2066 : AOI21_X1 port map( B1 => n809, B2 => n270, A => n811, ZN => n804);
   U2067 : XNOR2_X1 port map( A => n1920, B => n770, ZN => n695);
   U2068 : XNOR2_X1 port map( A => n904, B => n914, ZN => n206);
   U2069 : NOR2_X1 port map( A1 => n915, A2 => n907, ZN => n914);
   U2070 : AOI211_X1 port map( C1 => n1892, C2 => n910, A => n916, B => n917, 
                           ZN => n915);
   U2071 : XNOR2_X1 port map( A => n2143, B => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n560);
   U2072 : AOI21_X1 port map( B1 => n912, B2 => n911, A => n922, ZN => n917);
   U2073 : XNOR2_X1 port map( A => n924, B => n925, ZN => n217);
   U2074 : NAND2_X1 port map( A1 => n911, A2 => n2069, ZN => n924);
   U2075 : INV_X1 port map( A => n922, ZN => n2069);
   U2076 : OAI21_X1 port map( B1 => n2075, B2 => n2074, A => n2072, ZN => n886)
                           ;
   U2077 : OAI21_X1 port map( B1 => n2074, B2 => n2071, A => n2072, ZN => n885)
                           ;
   U2078 : INV_X1 port map( A => n159, ZN => n2095);
   U2079 : OAI21_X1 port map( B1 => n118, B2 => n1903, A => n2015, ZN => n124);
   U2080 : OAI21_X1 port map( B1 => n192, B2 => n1903, A => n2015, ZN => n194);
   U2081 : OAI21_X1 port map( B1 => n214, B2 => n1903, A => n2015, ZN => n216);
   U2082 : OAI21_X1 port map( B1 => n224, B2 => n1902, A => n2015, ZN => n226);
   U2083 : OAI21_X1 port map( B1 => n234, B2 => n1903, A => n2015, ZN => n236);
   U2084 : OAI21_X1 port map( B1 => n246, B2 => n1902, A => n2015, ZN => n248);
   U2085 : OAI21_X1 port map( B1 => n256, B2 => n1903, A => n2015, ZN => n258);
   U2086 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_2_port, A => n2015, 
                           ZN => n267);
   U2087 : OAI22_X1 port map( A1 => n1972, A2 => n1599, B1 => n1636, B2 => 
                           n1970, ZN => n1500);
   U2088 : OAI22_X1 port map( A1 => n1971, A2 => n1598, B1 => n1645, B2 => 
                           n1969, ZN => n1506);
   U2089 : OAI22_X1 port map( A1 => n1971, A2 => n1621, B1 => n1591, B2 => 
                           n1970, ZN => n1510);
   U2090 : NOR2_X1 port map( A1 => n916, A2 => n907, ZN => n905);
   U2091 : NOR2_X1 port map( A1 => n457, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, ZN => n732);
   U2092 : OAI22_X1 port map( A1 => n1974, A2 => n1593, B1 => n1707, B2 => 
                           n1970, ZN => n1484);
   U2093 : OAI22_X1 port map( A1 => n1634, A2 => n1963, B1 => n2035, B2 => 
                           n1961, ZN => n1567);
   U2094 : OAI22_X1 port map( A1 => n1635, A2 => n1963, B1 => n2034, B2 => 
                           n1961, ZN => n1566);
   U2095 : OAI22_X1 port map( A1 => n1637, A2 => n1963, B1 => n2033, B2 => 
                           n1961, ZN => n1565);
   U2096 : OAI21_X1 port map( B1 => n732, B2 => n2133, A => n733, ZN => n434);
   U2097 : OAI21_X1 port map( B1 => n729, B2 => n2098, A => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, ZN => n733);
   U2098 : OAI21_X1 port map( B1 => n2097, B2 => n2133, A => n728, ZN => n432);
   U2099 : OAI211_X1 port map( C1 => DATAPATH_IxThird_stxALU_IN1_29_port, C2 =>
                           n729, A => DATAPATH_IxThird_stxALU_IN1_28_port, B =>
                           n457, ZN => n728);
   U2100 : NOR2_X1 port map( A1 => n380, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, ZN => n377);
   U2101 : NOR2_X1 port map( A1 => n447, A2 => n1575, ZN => n443);
   U2102 : INV_X1 port map( A => CU_IxN24, ZN => n2001);
   U2103 : XNOR2_X1 port map( A => n244, B => n2083, ZN => n1291);
   U2104 : XNOR2_X1 port map( A => n814, B => n1774, ZN => 
                           DATAPATH_IxSecond_stxjump_target_3_port);
   U2105 : NAND2_X1 port map( A1 => n2087, A2 => n1677, ZN => n814);
   U2106 : INV_X1 port map( A => n1090, ZN => n2201);
   U2107 : OAI21_X1 port map( B1 => n2075, B2 => n900, A => n901, ZN => 
                           DATAPATH_IxSecond_stxjump_target_16_port);
   U2108 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_6_port, ZN => 
                           n2123);
   U2109 : NAND2_X1 port map( A1 => n695, A2 => n1794, ZN => n692);
   U2110 : NAND2_X1 port map( A1 => n650, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n648);
   U2111 : NAND2_X1 port map( A1 => n498, A2 => n1674, ZN => n492);
   U2112 : NAND2_X1 port map( A1 => n605, A2 => n1669, ZN => n600);
   U2113 : INV_X1 port map( A => n401, ZN => n2161);
   U2114 : NAND2_X1 port map( A1 => n388, A2 => n1791, ZN => n379);
   U2115 : OAI21_X1 port map( B1 => n783, B2 => n786, A => n600, ZN => n784);
   U2116 : NAND2_X1 port map( A1 => n601, A2 => n1655, ZN => n786);
   U2117 : INV_X1 port map( A => n913, ZN => n2070);
   U2118 : INV_X1 port map( A => n165, ZN => n2094);
   U2119 : AOI21_X1 port map( B1 => n2105, B2 => n2139, A => n507, ZN => n504);
   U2120 : INV_X1 port map( A => n495, ZN => n2139);
   U2121 : AND2_X1 port map( A1 => n2015, A2 => n289, ZN => n285);
   U2122 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_29_port, ZN => 
                           n2097);
   U2123 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_3_port, ZN => 
                           n2126);
   U2124 : OAI221_X1 port map( B1 => n2146, B2 => n607, C1 => n1912, C2 => n608
                           , A => n609, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_17_port);
   U2125 : AOI21_X1 port map( B1 => n1956, B2 => n1668, A => n1955, ZN => n607)
                           ;
   U2126 : XNOR2_X1 port map( A => n611, B => n2112, ZN => n608);
   U2127 : OAI21_X1 port map( B1 => n171, B2 => n1903, A => n2015, ZN => n169);
   U2128 : NAND2_X1 port map( A1 => n911, A2 => n912, ZN => n909);
   U2129 : NAND2_X1 port map( A1 => n380, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, ZN => n378);
   U2130 : NAND2_X1 port map( A1 => n447, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, ZN => n444);
   U2131 : OAI21_X1 port map( B1 => n748, B2 => n553, A => n540, ZN => n746);
   U2132 : BUF_X1 port map( A => n1939, Z => n1933);
   U2133 : BUF_X1 port map( A => n1939, Z => n1936);
   U2134 : BUF_X1 port map( A => n1939, Z => n1937);
   U2135 : BUF_X1 port map( A => n1939, Z => n1935);
   U2136 : BUF_X1 port map( A => n1939, Z => n1932);
   U2137 : BUF_X1 port map( A => n1939, Z => n1934);
   U2138 : BUF_X1 port map( A => n1864, Z => n1976);
   U2139 : BUF_X1 port map( A => n1864, Z => n1975);
   U2140 : BUF_X1 port map( A => n1864, Z => n1974);
   U2141 : BUF_X1 port map( A => n1864, Z => n1973);
   U2142 : BUF_X1 port map( A => n1864, Z => n1972);
   U2143 : BUF_X1 port map( A => n1864, Z => n1971);
   U2144 : INV_X1 port map( A => n877, ZN => n2075);
   U2145 : OAI21_X1 port map( B1 => n1634, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_12_port);
   U2146 : OAI21_X1 port map( B1 => n1635, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_13_port);
   U2147 : OAI21_X1 port map( B1 => n1637, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_14_port);
   U2148 : OAI21_X1 port map( B1 => n1646, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_29_port);
   U2149 : OAI21_X1 port map( B1 => n1386, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_31_port);
   U2150 : OAI21_X1 port map( B1 => n769, B2 => n336, A => n692, ZN => n767);
   U2151 : BUF_X1 port map( A => n1864, Z => n1977);
   U2152 : OAI21_X1 port map( B1 => n800, B2 => n801, A => n2198, ZN => n798);
   U2153 : BUF_X1 port map( A => n1939, Z => n1938);
   U2154 : BUF_X1 port map( A => n1689, Z => n1915);
   U2155 : NAND2_X1 port map( A1 => n1093, A2 => n1092, ZN => n1090);
   U2156 : INV_X1 port map( A => n878, ZN => n2071);
   U2157 : AOI21_X1 port map( B1 => n1956, B2 => n1655, A => n1955, ZN => n615)
                           ;
   U2158 : XNOR2_X1 port map( A => n2114, B => n619, ZN => n616);
   U2159 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_10_port, ZN => 
                           n2118);
   U2160 : INV_X1 port map( A => n1787, ZN => n2116);
   U2161 : INV_X1 port map( A => n171, ZN => n2203);
   U2162 : INV_X1 port map( A => n1138, ZN => n2042);
   U2163 : INV_X1 port map( A => n256, ZN => n2209);
   U2164 : INV_X1 port map( A => n246, ZN => n2208);
   U2165 : INV_X1 port map( A => n234, ZN => n2207);
   U2166 : INV_X1 port map( A => n224, ZN => n2206);
   U2167 : INV_X1 port map( A => n214, ZN => n2205);
   U2168 : INV_X1 port map( A => n192, ZN => n2204);
   U2169 : AND2_X1 port map( A1 => n730, A2 => n1783, ZN => n719);
   U2170 : INV_X1 port map( A => n789, ZN => n2135);
   U2171 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_26_port, ZN => 
                           n2103);
   U2172 : INV_X1 port map( A => n734, ZN => n2132);
   U2173 : INV_X1 port map( A => n770, ZN => n2154);
   U2174 : INV_X1 port map( A => n771, ZN => n2155);
   U2175 : INV_X1 port map( A => n894, ZN => n2074);
   U2176 : NAND2_X1 port map( A1 => n2072, A2 => n894, ZN => n874);
   U2177 : INV_X1 port map( A => n872, ZN => n2073);
   U2178 : INV_X1 port map( A => n91, ZN => n2005);
   U2179 : OAI21_X1 port map( B1 => CU_Ixcw_LUT_15_port, B2 => n1994, A => 
                           n1965, ZN => n91);
   U2180 : INV_X1 port map( A => n118, ZN => n2202);
   U2181 : INV_X1 port map( A => n735, ZN => n2134);
   U2182 : INV_X1 port map( A => n742, ZN => n2138);
   U2183 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_27_port, ZN => 
                           n2102);
   U2184 : INV_X1 port map( A => n271, ZN => n2084);
   U2185 : OR2_X1 port map( A1 => n730, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, ZN => n727);
   U2186 : AOI21_X1 port map( B1 => n597, B2 => n784, A => n585, ZN => n751);
   U2187 : NAND2_X1 port map( A1 => n2199, A2 => n809, ZN => n813);
   U2188 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_22_port, ZN => 
                           n2107);
   U2189 : INV_X1 port map( A => CU_IxN23, ZN => n2000);
   U2190 : INV_X1 port map( A => n811, ZN => n2199);
   U2191 : INV_X1 port map( A => n237, ZN => n2082);
   U2192 : INV_X1 port map( A => n47, ZN => n2058);
   U2193 : INV_X1 port map( A => n949, ZN => n2196);
   U2194 : OAI221_X1 port map( B1 => n1911, B2 => n572, C1 => n1889, C2 => n574
                           , A => n575, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_19_port);
   U2195 : INV_X1 port map( A => n1995, ZN => n1991);
   U2196 : NOR3_X1 port map( A1 => n2042, A2 => n1993, A3 => n2045, ZN => n28);
   U2197 : INV_X1 port map( A => n1982, ZN => n1981);
   U2198 : INV_X1 port map( A => n1865, ZN => n1956);
   U2199 : AOI21_X1 port map( B1 => n1639, B2 => n1915, A => n860, ZN => n851);
   U2200 : AOI21_X1 port map( B1 => n1640, B2 => n1916, A => n843, ZN => n834);
   U2201 : INV_X1 port map( A => n1865, ZN => n1957);
   U2202 : OAI21_X1 port map( B1 => n1929, B2 => n1605, A => n790, ZN => n421);
   U2203 : BUF_X1 port map( A => n334, Z => n1960);
   U2204 : NOR2_X1 port map( A1 => n605, A2 => n1669, ZN => n599);
   U2205 : NOR2_X1 port map( A1 => n695, A2 => n1794, ZN => n691);
   U2206 : NOR2_X1 port map( A1 => n498, A2 => n1674, ZN => n496);
   U2207 : NOR2_X1 port map( A1 => n650, A2 => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n646);
   U2208 : NOR2_X1 port map( A1 => n933, A2 => n941, ZN => n931);
   U2209 : OAI21_X1 port map( B1 => n949, B2 => n794, A => n950, ZN => n942);
   U2210 : OAI21_X1 port map( B1 => n690, B2 => n691, A => n692, ZN => n675);
   U2211 : NOR2_X1 port map( A1 => n1809, A2 => n337, ZN => n690);
   U2212 : NOR2_X1 port map( A1 => n569, A2 => n1786, ZN => n442);
   U2213 : OAI21_X1 port map( B1 => n598, B2 => n599, A => n600, ZN => n583);
   U2214 : NOR2_X1 port map( A1 => n1655, A2 => n601, ZN => n598);
   U2215 : OAI21_X1 port map( B1 => n545, B2 => n544, A => n540, ZN => n529);
   U2216 : NOR2_X1 port map( A1 => DATAPATH_IxThird_stxALU_IN1_20_port, A2 => 
                           n543, ZN => n545);
   U2217 : NOR2_X1 port map( A1 => n388, A2 => n1791, ZN => n376);
   U2218 : OAI21_X1 port map( B1 => n497, B2 => n496, A => n492, ZN => n480);
   U2219 : BUF_X1 port map( A => n334, Z => n1959);
   U2220 : BUF_X1 port map( A => n334, Z => n1958);
   U2221 : NOR2_X1 port map( A1 => n658, A2 => n1796, ZN => n649);
   U2222 : NAND2_X1 port map( A1 => n540, A2 => n541, ZN => n525);
   U2223 : INV_X1 port map( A => n544, ZN => n2108);
   U2224 : OAI21_X1 port map( B1 => n2127, B2 => n1865, A => n1603, ZN => n439)
                           ;
   U2225 : AOI21_X1 port map( B1 => n1916, B2 => n1638, A => n824, ZN => n821);
   U2226 : OAI21_X1 port map( B1 => n2126, B2 => n1865, A => n1603, ZN => n400)
                           ;
   U2227 : OAI21_X1 port map( B1 => n1917, B2 => n1638, A => n826, ZN => n825);
   U2228 : OAI21_X1 port map( B1 => n941, B2 => n942, A => n2195, ZN => n940);
   U2229 : BUF_X1 port map( A => n1916, Z => n1914);
   U2230 : INV_X1 port map( A => n418, ZN => n2159);
   U2231 : BUF_X1 port map( A => n1914, Z => n1917);
   U2232 : NAND2_X1 port map( A1 => n692, A2 => n693, ZN => n679);
   U2233 : INV_X1 port map( A => n691, ZN => n2119);
   U2234 : NAND2_X1 port map( A1 => n492, A2 => n493, ZN => n476);
   U2235 : INV_X1 port map( A => n496, ZN => n2104);
   U2236 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_16_port, ZN => 
                           n2113);
   U2237 : INV_X1 port map( A => n933, ZN => n2195);
   U2238 : INV_X1 port map( A => n805, ZN => n2198);
   U2239 : INV_X1 port map( A => n298, ZN => n2158);
   U2240 : INV_X1 port map( A => n705, ZN => n2129);
   U2241 : AOI21_X1 port map( B1 => n1786, B2 => n1956, A => n1955, ZN => n705)
                           ;
   U2242 : INV_X1 port map( A => n570, ZN => n2128);
   U2243 : AOI21_X1 port map( B1 => n1575, B2 => n1956, A => n1955, ZN => n570)
                           ;
   U2244 : INV_X1 port map( A => n292, ZN => n2096);
   U2245 : OAI221_X1 port map( B1 => n1860, B2 => n1615, C1 => n1431, C2 => 
                           n1951, A => n1050, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_12_port);
   U2246 : OAI221_X1 port map( B1 => n1860, B2 => n1604, C1 => n1436, C2 => 
                           n1950, A => n1007, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_17_port);
   U2247 : OAI221_X1 port map( B1 => n1871, B2 => n1593, C1 => n1434, C2 => 
                           n1951, A => n1046, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_15_port);
   U2248 : AOI211_X1 port map( C1 => n1637, C2 => n2076, A => n896, B => n1349,
                           ZN => n907);
   U2249 : NOR3_X1 port map( A1 => n2048, A2 => IRAM_DOUT(3), A3 => n2047, ZN 
                           => n1137);
   U2250 : NOR3_X1 port map( A1 => n1390, A2 => n1389, A3 => n1391, ZN => n256)
                           ;
   U2251 : NOR3_X1 port map( A1 => n1393, A2 => n1392, A3 => n2209, ZN => n246)
                           ;
   U2252 : NOR3_X1 port map( A1 => n1395, A2 => n1394, A3 => n2208, ZN => n234)
                           ;
   U2253 : NOR3_X1 port map( A1 => n1397, A2 => n1396, A3 => n2207, ZN => n224)
                           ;
   U2254 : NOR3_X1 port map( A1 => n1399, A2 => n1398, A3 => n2206, ZN => n214)
                           ;
   U2255 : NOR3_X1 port map( A1 => n1403, A2 => n1402, A3 => n198, ZN => n192);
   U2256 : AOI211_X1 port map( C1 => n2076, C2 => n1372, A => n896, B => n1350,
                           ZN => n878);
   U2257 : NOR2_X1 port map( A1 => n838, A2 => n839, ZN => n837);
   U2258 : AOI22_X1 port map( A1 => RF_WR_DATAx28x, A2 => n1943, B1 => 
                           RF_RD2_DATA(28), B2 => n1940, ZN => n1030);
   U2259 : AOI22_X1 port map( A1 => RF_WR_DATAx29x, A2 => n1943, B1 => 
                           RF_RD2_DATA(29), B2 => n1816, ZN => n1033);
   U2260 : OAI221_X1 port map( B1 => n1428, B2 => n1762, C1 => n1184, C2 => 
                           n1869, A => n1041, ZN => n770);
   U2261 : AOI22_X1 port map( A1 => RF_WR_DATAx9x, A2 => n1943, B1 => 
                           RF_RD2_DATA(9), B2 => n1940, ZN => n1041);
   U2262 : NAND2_X1 port map( A1 => n1205, A2 => n2093, ZN => n963);
   U2263 : NAND2_X1 port map( A1 => n1205, A2 => n2093, ZN => n1897);
   U2264 : NOR3_X1 port map( A1 => n1413, A2 => n1412, A3 => n132, ZN => n118);
   U2265 : AOI21_X1 port map( B1 => n1819, B2 => n1414, A => n124, ZN => n119);
   U2266 : OAI221_X1 port map( B1 => n1446, B2 => n1761, C1 => n1167, C2 => 
                           n1770, A => n1027, ZN => n789);
   U2267 : AOI22_X1 port map( A1 => RF_WR_DATAx27x, A2 => n1943, B1 => 
                           RF_RD2_DATA(27), B2 => n1940, ZN => n1027);
   U2268 : AOI22_X1 port map( A1 => n2083, A2 => n2197, B1 => n1384, B2 => 
                           n1343, ZN => n792);
   U2269 : INV_X1 port map( A => n794, ZN => n2197);
   U2270 : XNOR2_X1 port map( A => n1364, B => n1386, ZN => n829);
   U2271 : NAND4_X1 port map( A1 => IRAM_DOUT(2), A2 => IRAM_DOUT(6), A3 => 
                           IRAM_DOUT(3), A4 => n1141, ZN => n1134);
   U2272 : NOR4_X1 port map( A1 => IRAM_DOUT(4), A2 => n2048, A3 => n2047, A4 
                           => n2044, ZN => n1141);
   U2273 : AOI211_X1 port map( C1 => n2076, C2 => n1374, A => n896, B => n1352,
                           ZN => n872);
   U2274 : OAI21_X1 port map( B1 => n1140, B2 => n2042, A => n1134, ZN => 
                           CU_IxN23);
   U2275 : AOI22_X1 port map( A1 => n27, A2 => n2045, B1 => IRAM_DOUT(4), B2 =>
                           n2044, ZN => n1140);
   U2276 : NOR4_X1 port map( A1 => n1417, A2 => n1902, A3 => n101, A4 => 
                           IRAM_ADD_31_port, ZN => n99);
   U2277 : NOR4_X1 port map( A1 => n1412, A2 => n132, A3 => n1901, A4 => 
                           IRAM_ADD_26_port, ZN => n137);
   U2278 : NOR4_X1 port map( A1 => n1406, A2 => n172, A3 => n1901, A4 => 
                           IRAM_ADD_20_port, ZN => n177);
   U2279 : NOR4_X1 port map( A1 => n1402, A2 => n198, A3 => n1901, A4 => 
                           IRAM_ADD_16_port, ZN => n203);
   U2280 : AOI21_X1 port map( B1 => n1819, B2 => n1390, A => n267, ZN => n266);
   U2281 : OAI222_X1 port map( A1 => n1213, A2 => n1907, B1 => n1387, B2 => 
                           n285, C1 => n1338, C2 => n1905, ZN => n1547);
   U2282 : OAI222_X1 port map( A1 => n1905, A2 => n49, B1 => n1388, B2 => n285,
                           C1 => n1214, C2 => n1907, ZN => n1546);
   U2283 : NOR2_X1 port map( A1 => n2044, A2 => IRAM_DOUT(2), ZN => n27);
   U2284 : NOR3_X1 port map( A1 => n1407, A2 => n1406, A3 => n172, ZN => n171);
   U2285 : AOI22_X1 port map( A1 => RF_WR_DATAx11x, A2 => n1578, B1 => 
                           RF_RD2_DATA(11), B2 => n985, ZN => n1059);
   U2286 : OAI21_X1 port map( B1 => n1765, B2 => n1241, A => n1677, ZN => n280)
                           ;
   U2287 : INV_X1 port map( A => n1051, ZN => n2152);
   U2288 : OAI221_X1 port map( B1 => n1431, B2 => n1761, C1 => n1182, C2 => 
                           n1869, A => n1052, ZN => n1051);
   U2289 : AOI22_X1 port map( A1 => RF_WR_DATAx12x, A2 => n1577, B1 => 
                           RF_RD2_DATA(12), B2 => n985, ZN => n1052);
   U2290 : OAI221_X1 port map( B1 => n1443, B2 => n1762, C1 => n1172, C2 => 
                           n1868, A => n1020, ZN => n742);
   U2291 : OAI221_X1 port map( B1 => n1439, B2 => n1762, C1 => n1178, C2 => 
                           n1869, A => n995, ZN => n750);
   U2292 : OAI221_X1 port map( B1 => n1860, B2 => n1596, C1 => n1433, C2 => 
                           n1951, A => n1043, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_14_port);
   U2293 : OAI221_X1 port map( B1 => n1861, B2 => n1606, C1 => n1428, C2 => 
                           n1951, A => n1040, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_9_port);
   U2294 : NOR2_X1 port map( A1 => n1197, A2 => n1298, ZN => n298);
   U2295 : AOI21_X1 port map( B1 => n113, B2 => IRAM_ADD_29_port, A => n115, ZN
                           => n112);
   U2296 : NOR3_X1 port map( A1 => IRAM_ADD_29_port, A2 => n110, A3 => n1901, 
                           ZN => n115);
   U2297 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_28_port, A => n119, 
                           ZN => n113);
   U2298 : NOR2_X1 port map( A1 => n1341, A2 => n1381, ZN => n811);
   U2299 : AOI21_X1 port map( B1 => n2076, B2 => n1371, A => n896, ZN => n913);
   U2300 : XNOR2_X1 port map( A => n2079, B => n1346, ZN => n930);
   U2301 : NAND4_X1 port map( A1 => IRAM_DOUT(6), A2 => n27, A3 => n1137, A4 =>
                           n2045, ZN => n26);
   U2302 : OAI221_X1 port map( B1 => n1904, B2 => n47, C1 => n1234, C2 => n1906
                           , A => n120, ZN => n1519);
   U2303 : AOI21_X1 port map( B1 => n2006, B2 => IRAM_ADD_28_port, A => n122, 
                           ZN => n120);
   U2304 : NOR4_X1 port map( A1 => n1414, A2 => n2202, A3 => n1901, A4 => 
                           IRAM_ADD_28_port, ZN => n122);
   U2305 : INV_X1 port map( A => n119, ZN => n2006);
   U2306 : OAI221_X1 port map( B1 => n1904, B2 => n2062, C1 => n1226, C2 => 
                           n1906, A => n174, ZN => n1527);
   U2307 : AOI21_X1 port map( B1 => n175, B2 => IRAM_ADD_20_port, A => n177, ZN
                           => n174);
   U2308 : INV_X1 port map( A => n1292, ZN => n2062);
   U2309 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_19_port, A => n179, 
                           ZN => n175);
   U2310 : OAI221_X1 port map( B1 => n1231, B2 => n1906, C1 => n1773, C2 => 
                           n1904, A => n141, ZN => n1522);
   U2311 : AOI21_X1 port map( B1 => n2011, B2 => IRAM_ADD_25_port, A => n143, 
                           ZN => n141);
   U2312 : INV_X1 port map( A => n139, ZN => n2011);
   U2313 : OAI221_X1 port map( B1 => n1237, B2 => n1907, C1 => n2059, C2 => 
                           n1905, A => n96, ZN => n1516);
   U2314 : AOI21_X1 port map( B1 => n97, B2 => IRAM_ADD_31_port, A => n99, ZN 
                           => n96);
   U2315 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_31_port, ZN 
                           => n2059);
   U2316 : OAI21_X1 port map( B1 => n1902, B2 => IRAM_ADD_30_port, A => n103, 
                           ZN => n97);
   U2317 : OAI221_X1 port map( B1 => n1236, B2 => n1906, C1 => n2060, C2 => 
                           n1904, A => n105, ZN => n1517);
   U2318 : AOI22_X1 port map( A1 => n106, A2 => n1417, B1 => n2012, B2 => 
                           IRAM_ADD_30_port, ZN => n105);
   U2319 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_30_port, ZN 
                           => n2060);
   U2320 : NOR2_X1 port map( A1 => n1903, A2 => n101, ZN => n106);
   U2321 : OAI221_X1 port map( B1 => n1904, B2 => n46, C1 => n1230, C2 => n1906
                           , A => n145, ZN => n1523);
   U2322 : AOI21_X1 port map( B1 => n146, B2 => IRAM_ADD_24_port, A => n148, ZN
                           => n145);
   U2323 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_23_port, A => n150, 
                           ZN => n146);
   U2324 : NOR4_X1 port map( A1 => n1410, A2 => n144, A3 => n1901, A4 => 
                           IRAM_ADD_24_port, ZN => n148);
   U2325 : OAI221_X1 port map( B1 => n1233, B2 => n1906, C1 => n2055, C2 => 
                           n1904, A => n129, ZN => n1520);
   U2326 : AOI21_X1 port map( B1 => n124, B2 => IRAM_ADD_27_port, A => n130, ZN
                           => n129);
   U2327 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_27_port, ZN 
                           => n2055);
   U2328 : NOR3_X1 port map( A1 => IRAM_ADD_27_port, A2 => n2202, A3 => n1901, 
                           ZN => n130);
   U2329 : OAI221_X1 port map( B1 => n1232, B2 => n1906, C1 => n2056, C2 => 
                           n1904, A => n134, ZN => n1521);
   U2330 : AOI21_X1 port map( B1 => n135, B2 => IRAM_ADD_26_port, A => n137, ZN
                           => n134);
   U2331 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_26_port, ZN 
                           => n2056);
   U2332 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_25_port, A => n139, 
                           ZN => n135);
   U2333 : OAI221_X1 port map( B1 => n1227, B2 => n1906, C1 => n2052, C2 => 
                           n1904, A => n167, ZN => n1526);
   U2334 : AOI22_X1 port map( A1 => n168, A2 => n1408, B1 => n169, B2 => 
                           IRAM_ADD_21_port, ZN => n167);
   U2335 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_21_port, ZN 
                           => n2052);
   U2336 : OAI221_X1 port map( B1 => n1229, B2 => n1906, C1 => n2051, C2 => 
                           n1904, A => n154, ZN => n1524);
   U2337 : AOI21_X1 port map( B1 => n2010, B2 => IRAM_ADD_23_port, A => n156, 
                           ZN => n154);
   U2338 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_23_port, ZN 
                           => n2051);
   U2339 : INV_X1 port map( A => n150, ZN => n2010);
   U2340 : OAI221_X1 port map( B1 => n1224, B2 => n1907, C1 => n2064, C2 => 
                           n1904, A => n196, ZN => n1530);
   U2341 : AOI21_X1 port map( B1 => n194, B2 => IRAM_ADD_17_port, A => n197, ZN
                           => n196);
   U2342 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_17_port, ZN 
                           => n2064);
   U2343 : NOR3_X1 port map( A1 => IRAM_ADD_17_port, A2 => n2204, A3 => n1902, 
                           ZN => n197);
   U2344 : OAI221_X1 port map( B1 => n1219, B2 => n1907, C1 => n1905, C2 => 
                           n237, A => n238, ZN => n1538);
   U2345 : AOI21_X1 port map( B1 => n236, B2 => IRAM_ADD_9_port, A => n239, ZN 
                           => n238);
   U2346 : NOR3_X1 port map( A1 => IRAM_ADD_9_port, A2 => n2207, A3 => n1902, 
                           ZN => n239);
   U2347 : OAI221_X1 port map( B1 => n1217, B2 => n1907, C1 => n2081, C2 => 
                           n1905, A => n260, ZN => n1542);
   U2348 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_5_port, ZN =>
                           n2081);
   U2349 : AOI21_X1 port map( B1 => n258, B2 => IRAM_ADD_5_port, A => n261, ZN 
                           => n260);
   U2350 : NOR3_X1 port map( A1 => IRAM_ADD_5_port, A2 => n2209, A3 => n1901, 
                           ZN => n261);
   U2351 : OAI221_X1 port map( B1 => n1904, B2 => n48, C1 => n1216, C2 => n1906
                           , A => n262, ZN => n1543);
   U2352 : AOI21_X1 port map( B1 => n2007, B2 => IRAM_ADD_4_port, A => n265, ZN
                           => n262);
   U2353 : NOR4_X1 port map( A1 => n1389, A2 => n1390, A3 => n1901, A4 => 
                           IRAM_ADD_4_port, ZN => n265);
   U2354 : INV_X1 port map( A => n266, ZN => n2007);
   U2355 : OAI221_X1 port map( B1 => n1215, B2 => n1907, C1 => n2086, C2 => 
                           n1905, A => n273, ZN => n1544);
   U2356 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_3_port, ZN =>
                           n2086);
   U2357 : AOI21_X1 port map( B1 => n267, B2 => IRAM_ADD_3_port, A => n275, ZN 
                           => n273);
   U2358 : NOR3_X1 port map( A1 => IRAM_ADD_3_port, A2 => n1389, A3 => n1901, 
                           ZN => n275);
   U2359 : OAI221_X1 port map( B1 => n1225, B2 => n1906, C1 => n1905, C2 => 
                           n182, A => n183, ZN => n1528);
   U2360 : AOI21_X1 port map( B1 => n2009, B2 => IRAM_ADD_19_port, A => n185, 
                           ZN => n183);
   U2361 : INV_X1 port map( A => n179, ZN => n2009);
   U2362 : NOR3_X1 port map( A1 => IRAM_ADD_19_port, A2 => n172, A3 => n1902, 
                           ZN => n185);
   U2363 : OAI221_X1 port map( B1 => n1223, B2 => n1907, C1 => n2063, C2 => 
                           n1905, A => n200, ZN => n1531);
   U2364 : AOI21_X1 port map( B1 => n201, B2 => IRAM_ADD_16_port, A => n203, ZN
                           => n200);
   U2365 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_16_port, ZN 
                           => n2063);
   U2366 : OAI21_X1 port map( B1 => n1903, B2 => IRAM_ADD_15_port, A => n205, 
                           ZN => n201);
   U2367 : OAI221_X1 port map( B1 => n1222, B2 => n1907, C1 => n1905, C2 => 
                           n206, A => n207, ZN => n1532);
   U2368 : AOI21_X1 port map( B1 => n2008, B2 => IRAM_ADD_15_port, A => n209, 
                           ZN => n207);
   U2369 : INV_X1 port map( A => n205, ZN => n2008);
   U2370 : NOR3_X1 port map( A1 => IRAM_ADD_15_port, A2 => n198, A3 => n1902, 
                           ZN => n209);
   U2371 : OAI221_X1 port map( B1 => n1221, B2 => n1907, C1 => n217, C2 => 
                           n1905, A => n218, ZN => n1534);
   U2372 : AOI21_X1 port map( B1 => n216, B2 => IRAM_ADD_13_port, A => n219, ZN
                           => n218);
   U2373 : NOR3_X1 port map( A1 => IRAM_ADD_13_port, A2 => n2205, A3 => n1902, 
                           ZN => n219);
   U2374 : OAI221_X1 port map( B1 => n1901, B2 => IRAM_ADD_2_port, C1 => n1905,
                           C2 => n2088, A => n278, ZN => n1545);
   U2375 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_2_port, B1 => n109, 
                           B2 => IRAM_ADD_2_port, ZN => n278);
   U2376 : INV_X1 port map( A => n1296, ZN => n2088);
   U2377 : INV_X1 port map( A => n1076, ZN => RF_WR_DATAx5x);
   U2378 : OAI22_X1 port map( A1 => n1932, A2 => DATAPATH_IxLMD_DATA_5_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_5_port, ZN 
                           => n1076);
   U2379 : NOR2_X1 port map( A1 => n1408, A2 => n2203, ZN => n164);
   U2380 : XNOR2_X1 port map( A => n913, B => n1257, ZN => n904);
   U2381 : INV_X1 port map( A => n1031, ZN => RF_WR_DATAx28x);
   U2382 : OAI22_X1 port map( A1 => n1935, A2 => DATAPATH_IxLMD_DATA_28_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_28_port, 
                           ZN => n1031);
   U2383 : NOR2_X1 port map( A1 => n1343, A2 => n1384, ZN => n794);
   U2384 : XNOR2_X1 port map( A => n1363, B => n1386, ZN => n830);
   U2385 : NOR2_X1 port map( A1 => n854, A2 => n855, ZN => n853);
   U2386 : XNOR2_X1 port map( A => n1163, B => n1146, ZN => n1102);
   U2387 : AOI21_X1 port map( B1 => n294, B2 => n298, A => n1197, ZN => n326);
   U2388 : NOR3_X1 port map( A1 => IRAM_ADD_25_port, A2 => n132, A3 => n1901, 
                           ZN => n143);
   U2389 : OAI221_X1 port map( B1 => n1220, B2 => n1907, C1 => n2078, C2 => 
                           n1905, A => n228, ZN => n1536);
   U2390 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_11_port, ZN 
                           => n2078);
   U2391 : AOI21_X1 port map( B1 => n226, B2 => IRAM_ADD_11_port, A => n229, ZN
                           => n228);
   U2392 : NOR3_X1 port map( A1 => IRAM_ADD_11_port, A2 => n2206, A3 => n1902, 
                           ZN => n229);
   U2393 : OAI221_X1 port map( B1 => n1218, B2 => n1907, C1 => n2080, C2 => 
                           n1905, A => n250, ZN => n1540);
   U2394 : INV_X1 port map( A => DATAPATH_IxSecond_stxjump_target_7_port, ZN =>
                           n2080);
   U2395 : AOI21_X1 port map( B1 => n248, B2 => IRAM_ADD_7_port, A => n251, ZN 
                           => n250);
   U2396 : NOR3_X1 port map( A1 => IRAM_ADD_7_port, A2 => n2208, A3 => n1902, 
                           ZN => n251);
   U2397 : INV_X1 port map( A => CU_Ixcw_LUT_16_port, ZN => n2041);
   U2398 : OAI22_X1 port map( A1 => n1975, A2 => n1612, B1 => n1354, B2 => 
                           n1969, ZN => n1474);
   U2399 : OAI22_X1 port map( A1 => n1376, A2 => n961, B1 => n1366, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_0_port);
   U2400 : OAI22_X1 port map( A1 => n1377, A2 => n961, B1 => n1367, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_1_port);
   U2401 : OAI22_X1 port map( A1 => n1378, A2 => n961, B1 => n1368, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_2_port);
   U2402 : OAI22_X1 port map( A1 => n1379, A2 => n961, B1 => n1369, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_3_port);
   U2403 : OAI22_X1 port map( A1 => n1380, A2 => n961, B1 => n1370, B2 => n962,
                           ZN => DATAPATH_IxSecond_stximm_extended_4_port);
   U2404 : OAI22_X1 port map( A1 => n1976, A2 => n1608, B1 => n1362, B2 => 
                           n1969, ZN => n1458);
   U2405 : OAI22_X1 port map( A1 => n1975, A2 => n1595, B1 => n1358, B2 => 
                           n1969, ZN => n1466);
   U2406 : OAI22_X1 port map( A1 => n1972, A2 => n1594, B1 => n1343, B2 => 
                           n1970, ZN => n1498);
   U2407 : OAI22_X1 port map( A1 => n1972, A2 => n1606, B1 => n1344, B2 => 
                           n1970, ZN => n1496);
   U2408 : XNOR2_X1 port map( A => n867, B => n1353, ZN => n869);
   U2409 : OAI22_X1 port map( A1 => n1976, A2 => n1607, B1 => n1363, B2 => 
                           n1969, ZN => n1456);
   U2410 : OAI22_X1 port map( A1 => n1976, A2 => n1613, B1 => n1359, B2 => 
                           n1969, ZN => n1464);
   U2411 : OAI22_X1 port map( A1 => n1975, A2 => n1618, B1 => n1355, B2 => 
                           n1969, ZN => n1472);
   U2412 : OAI22_X1 port map( A1 => n1900, A2 => n1591, B1 => n1389, B2 => 
                           n1968, ZN => n1511);
   U2413 : OAI22_X1 port map( A1 => n1355, A2 => n1899, B1 => n1408, B2 => 
                           n1966, ZN => n1473);
   U2414 : OAI22_X1 port map( A1 => n1340, A2 => n1898, B1 => n1390, B2 => 
                           n1968, ZN => n1509);
   U2415 : OAI221_X1 port map( B1 => n1445, B2 => n1762, C1 => n1168, C2 => 
                           n1769, A => n1024, ZN => n488);
   U2416 : AOI22_X1 port map( A1 => RF_WR_DATAx26x, A2 => n1943, B1 => 
                           RF_RD2_DATA(26), B2 => n1940, ZN => n1024);
   U2417 : OAI221_X1 port map( B1 => n1427, B2 => n1761, C1 => n1185, C2 => 
                           n1868, A => n1038, ZN => n771);
   U2418 : AOI22_X1 port map( A1 => RF_WR_DATAx8x, A2 => n1943, B1 => 
                           RF_RD2_DATA(8), B2 => n985, ZN => n1038);
   U2419 : OAI22_X1 port map( A1 => n1972, A2 => n1620, B1 => n1342, B2 => 
                           n1969, ZN => n1502);
   U2420 : OAI22_X1 port map( A1 => n1972, A2 => n1609, B1 => n1341, B2 => 
                           n1969, ZN => n1504);
   U2421 : OAI22_X1 port map( A1 => n1971, A2 => n1619, B1 => n1340, B2 => 
                           n1970, ZN => n1508);
   U2422 : OAI22_X1 port map( A1 => n1971, A2 => n1625, B1 => n1338, B2 => 
                           n1969, ZN => n1514);
   U2423 : OAI22_X1 port map( A1 => n1971, A2 => n1610, B1 => n1339, B2 => 
                           n1970, ZN => n1512);
   U2424 : OAI22_X1 port map( A1 => n1409, A2 => n2015, B1 => n109, B2 => n158,
                           ZN => n1525);
   U2425 : AOI211_X1 port map( C1 => n159, C2 => 
                           DATAPATH_IxSecond_stxjump_target_22_port, A => n160,
                           B => n161, ZN => n158);
   U2426 : OAI21_X1 port map( B1 => n1228, B2 => n165, A => n1991, ZN => n160);
   U2427 : NOR3_X1 port map( A1 => n162, A2 => n2094, A3 => n159, ZN => n161);
   U2428 : OAI22_X1 port map( A1 => n1974, A2 => n1600, B1 => n1353, B2 => 
                           n1970, ZN => n1476);
   U2429 : OAI22_X1 port map( A1 => n1973, A2 => n1626, B1 => n1346, B2 => 
                           n1970, ZN => n1492);
   U2430 : OAI22_X1 port map( A1 => n1977, A2 => n1616, B1 => n1364, B2 => 
                           n1969, ZN => n1454);
   U2431 : OAI22_X1 port map( A1 => n1976, A2 => n1627, B1 => n1360, B2 => 
                           n1969, ZN => n1462);
   U2432 : OAI22_X1 port map( A1 => n1975, A2 => n1614, B1 => n1356, B2 => 
                           n1969, ZN => n1470);
   U2433 : OAI22_X1 port map( A1 => n1346, A2 => n1898, B1 => n1398, B2 => 
                           n1967, ZN => n1493);
   U2434 : OAI22_X1 port map( A1 => n1344, A2 => n1898, B1 => n1396, B2 => 
                           n1967, ZN => n1497);
   U2435 : OAI22_X1 port map( A1 => n1900, A2 => n1636, B1 => n1394, B2 => 
                           n1968, ZN => n1501);
   U2436 : OAI22_X1 port map( A1 => n1341, A2 => n1898, B1 => n1392, B2 => 
                           n1968, ZN => n1505);
   U2437 : OAI221_X1 port map( B1 => n1880, B2 => n1595, C1 => n1443, C2 => 
                           n1950, A => n1019, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_24_port);
   U2438 : OAI22_X1 port map( A1 => n1973, A2 => n1596, B1 => n1349, B2 => 
                           n1970, ZN => n1486);
   U2439 : OAI22_X1 port map( A1 => n1351, A2 => n1899, B1 => n1404, B2 => 
                           n1967, ZN => n1481);
   U2440 : OAI22_X1 port map( A1 => n1348, A2 => n1898, B1 => n1400, B2 => 
                           n1967, ZN => n1489);
   U2441 : OAI22_X1 port map( A1 => n1353, A2 => n1899, B1 => n1406, B2 => 
                           n1967, ZN => n1477);
   U2442 : OAI22_X1 port map( A1 => n1900, A2 => n1707, B1 => n1402, B2 => 
                           n1967, ZN => n1485);
   U2443 : OAI22_X1 port map( A1 => n1357, A2 => n1899, B1 => n1410, B2 => 
                           n1966, ZN => n1469);
   U2444 : OAI22_X1 port map( A1 => n1361, A2 => n1900, B1 => n1414, B2 => 
                           n1966, ZN => n1461);
   U2445 : OAI22_X1 port map( A1 => n1347, A2 => n1898, B1 => n1399, B2 => 
                           n1967, ZN => n1491);
   U2446 : OAI22_X1 port map( A1 => n1345, A2 => n1898, B1 => n1397, B2 => 
                           n1967, ZN => n1495);
   U2447 : OAI22_X1 port map( A1 => n1343, A2 => n1898, B1 => n1395, B2 => 
                           n1967, ZN => n1499);
   U2448 : OAI22_X1 port map( A1 => n1342, A2 => n1898, B1 => n1393, B2 => 
                           n1968, ZN => n1503);
   U2449 : OAI22_X1 port map( A1 => n1352, A2 => n1899, B1 => n1405, B2 => 
                           n1967, ZN => n1479);
   U2450 : OAI22_X1 port map( A1 => n1349, A2 => n1898, B1 => n1401, B2 => 
                           n1967, ZN => n1487);
   U2451 : OAI22_X1 port map( A1 => n1976, A2 => n1628, B1 => n1361, B2 => 
                           n1969, ZN => n1460);
   U2452 : OAI22_X1 port map( A1 => n1975, A2 => n1617, B1 => n1357, B2 => 
                           n1969, ZN => n1468);
   U2453 : OAI22_X1 port map( A1 => n1356, A2 => n1899, B1 => n1409, B2 => 
                           n1966, ZN => n1471);
   U2454 : OAI22_X1 port map( A1 => n1973, A2 => n1629, B1 => n1345, B2 => 
                           n1970, ZN => n1494);
   U2455 : OAI22_X1 port map( A1 => n1974, A2 => n1611, B1 => n1352, B2 => 
                           n1970, ZN => n1478);
   U2456 : OAI22_X1 port map( A1 => n1974, A2 => n1604, B1 => n1351, B2 => 
                           n1970, ZN => n1480);
   U2457 : OAI22_X1 port map( A1 => n1974, A2 => n1597, B1 => n1350, B2 => 
                           n1970, ZN => n1482);
   U2458 : OAI22_X1 port map( A1 => n1973, A2 => n1630, B1 => n1348, B2 => 
                           n1970, ZN => n1488);
   U2459 : OAI22_X1 port map( A1 => n1973, A2 => n1615, B1 => n1347, B2 => 
                           n1970, ZN => n1490);
   U2460 : OAI22_X1 port map( A1 => n1900, A2 => n1645, B1 => n1391, B2 => 
                           n1968, ZN => n1507);
   U2461 : OAI22_X1 port map( A1 => n1338, A2 => n1898, B1 => n1387, B2 => 
                           n1968, ZN => n1515);
   U2462 : OAI22_X1 port map( A1 => n1339, A2 => n1898, B1 => n1388, B2 => 
                           n1968, ZN => n1513);
   U2463 : OAI22_X1 port map( A1 => n1977, A2 => n1622, B1 => n1365, B2 => 
                           n1969, ZN => n1452);
   U2464 : OAI22_X1 port map( A1 => n1359, A2 => n1899, B1 => n1412, B2 => 
                           n1966, ZN => n1465);
   U2465 : OAI22_X1 port map( A1 => n1360, A2 => n1899, B1 => n1413, B2 => 
                           n1966, ZN => n1463);
   U2466 : OAI22_X1 port map( A1 => n1354, A2 => n1899, B1 => n1407, B2 => 
                           n1966, ZN => n1475);
   U2467 : OAI22_X1 port map( A1 => n1350, A2 => n1899, B1 => n1403, B2 => 
                           n1967, ZN => n1483);
   U2468 : OAI22_X1 port map( A1 => n1358, A2 => n1899, B1 => n1411, B2 => 
                           n1966, ZN => n1467);
   U2469 : OAI22_X1 port map( A1 => n1364, A2 => n1900, B1 => n1417, B2 => 
                           n1966, ZN => n1455);
   U2470 : NOR2_X1 port map( A1 => n956, A2 => n1244, ZN => n271);
   U2471 : OAI22_X1 port map( A1 => n1366, A2 => n1963, B1 => n1961, B2 => 
                           n2040, ZN => n1572);
   U2472 : INV_X1 port map( A => IRAM_DOUT(7), ZN => n2040);
   U2473 : OAI22_X1 port map( A1 => n1367, A2 => n1963, B1 => n1962, B2 => 
                           n2039, ZN => n1571);
   U2474 : INV_X1 port map( A => IRAM_DOUT(8), ZN => n2039);
   U2475 : OAI22_X1 port map( A1 => n1368, A2 => n1963, B1 => n1962, B2 => 
                           n2038, ZN => n1570);
   U2476 : INV_X1 port map( A => IRAM_DOUT(9), ZN => n2038);
   U2477 : OAI22_X1 port map( A1 => n1369, A2 => n1963, B1 => n1962, B2 => 
                           n2037, ZN => n1569);
   U2478 : INV_X1 port map( A => IRAM_DOUT(10), ZN => n2037);
   U2479 : OAI22_X1 port map( A1 => n1370, A2 => n1963, B1 => n1962, B2 => 
                           n2036, ZN => n1568);
   U2480 : INV_X1 port map( A => IRAM_DOUT(11), ZN => n2036);
   U2481 : OAI22_X1 port map( A1 => n1371, A2 => n1963, B1 => n1962, B2 => 
                           n2032, ZN => n1564);
   U2482 : INV_X1 port map( A => IRAM_DOUT(15), ZN => n2032);
   U2483 : OAI22_X1 port map( A1 => n1372, A2 => n1963, B1 => n1962, B2 => 
                           n2031, ZN => n1563);
   U2484 : INV_X1 port map( A => IRAM_DOUT(16), ZN => n2031);
   U2485 : OAI22_X1 port map( A1 => n1373, A2 => n1963, B1 => n1962, B2 => 
                           n2030, ZN => n1562);
   U2486 : INV_X1 port map( A => IRAM_DOUT(17), ZN => n2030);
   U2487 : OAI22_X1 port map( A1 => n1374, A2 => n1964, B1 => n1962, B2 => 
                           n2029, ZN => n1561);
   U2488 : INV_X1 port map( A => IRAM_DOUT(18), ZN => n2029);
   U2489 : OAI22_X1 port map( A1 => n1375, A2 => n1964, B1 => n1962, B2 => 
                           n2028, ZN => n1560);
   U2490 : INV_X1 port map( A => IRAM_DOUT(19), ZN => n2028);
   U2491 : OAI22_X1 port map( A1 => n1376, A2 => n1964, B1 => n1962, B2 => 
                           n2027, ZN => n1559);
   U2492 : INV_X1 port map( A => IRAM_DOUT(20), ZN => n2027);
   U2493 : OAI22_X1 port map( A1 => n1377, A2 => n1964, B1 => n1962, B2 => 
                           n2026, ZN => n1558);
   U2494 : INV_X1 port map( A => IRAM_DOUT(21), ZN => n2026);
   U2495 : OAI22_X1 port map( A1 => n1378, A2 => n1964, B1 => n1962, B2 => 
                           n2025, ZN => n1557);
   U2496 : INV_X1 port map( A => IRAM_DOUT(22), ZN => n2025);
   U2497 : OAI22_X1 port map( A1 => n1379, A2 => n1964, B1 => n1961, B2 => 
                           n2024, ZN => n1556);
   U2498 : INV_X1 port map( A => IRAM_DOUT(23), ZN => n2024);
   U2499 : OAI22_X1 port map( A1 => n1380, A2 => n1964, B1 => n1961, B2 => 
                           n2023, ZN => n1555);
   U2500 : INV_X1 port map( A => IRAM_DOUT(24), ZN => n2023);
   U2501 : OAI22_X1 port map( A1 => n1381, A2 => n1964, B1 => n1961, B2 => 
                           n2022, ZN => n1554);
   U2502 : INV_X1 port map( A => IRAM_DOUT(25), ZN => n2022);
   U2503 : OAI22_X1 port map( A1 => n1382, A2 => n1964, B1 => n1961, B2 => 
                           n2021, ZN => n1553);
   U2504 : INV_X1 port map( A => IRAM_DOUT(26), ZN => n2021);
   U2505 : OAI22_X1 port map( A1 => n1383, A2 => n1964, B1 => n1961, B2 => 
                           n2020, ZN => n1552);
   U2506 : INV_X1 port map( A => IRAM_DOUT(27), ZN => n2020);
   U2507 : OAI22_X1 port map( A1 => n1384, A2 => n1964, B1 => n1961, B2 => 
                           n2019, ZN => n1551);
   U2508 : INV_X1 port map( A => IRAM_DOUT(28), ZN => n2019);
   U2509 : OAI22_X1 port map( A1 => n1646, A2 => n1964, B1 => n1961, B2 => 
                           n2018, ZN => n1550);
   U2510 : INV_X1 port map( A => IRAM_DOUT(29), ZN => n2018);
   U2511 : OAI22_X1 port map( A1 => n1385, A2 => n1965, B1 => n1961, B2 => 
                           n2017, ZN => n1549);
   U2512 : INV_X1 port map( A => IRAM_DOUT(30), ZN => n2017);
   U2513 : OAI22_X1 port map( A1 => n1386, A2 => n1965, B1 => n1962, B2 => 
                           n2016, ZN => n1548);
   U2514 : INV_X1 port map( A => IRAM_DOUT(31), ZN => n2016);
   U2515 : OAI22_X1 port map( A1 => n1365, A2 => n1899, B1 => n1418, B2 => 
                           n1966, ZN => n1453);
   U2516 : OAI22_X1 port map( A1 => n1363, A2 => n1900, B1 => n1416, B2 => 
                           n1966, ZN => n1457);
   U2517 : OAI22_X1 port map( A1 => n1362, A2 => n1900, B1 => n1415, B2 => 
                           n1966, ZN => n1459);
   U2518 : NOR2_X1 port map( A1 => n1646, A2 => n1344, ZN => n949);
   U2519 : NOR2_X1 port map( A1 => n2046, A2 => IRAM_DOUT(6), ZN => n1138);
   U2520 : INV_X1 port map( A => n1137, ZN => n2046);
   U2521 : XNOR2_X1 port map( A => n865, B => n852, ZN => 
                           DATAPATH_IxSecond_stxjump_target_21_port);
   U2522 : OAI21_X1 port map( B1 => n2053, B2 => n1386, A => n1354, ZN => n866)
                           ;
   U2523 : XNOR2_X1 port map( A => n1344, B => n1646, ZN => n791);
   U2524 : XNOR2_X1 port map( A => n1576, B => n836, ZN => 
                           DATAPATH_IxSecond_stxjump_target_25_port);
   U2525 : NOR2_X1 port map( A1 => n1382, A2 => n1342, ZN => n805);
   U2526 : AOI22_X1 port map( A1 => RF_WR_DATAx14x, A2 => n1943, B1 => 
                           RF_RD2_DATA(14), B2 => n985, ZN => n1044);
   U2527 : INV_X1 port map( A => IRAM_DOUT(4), ZN => n2045);
   U2528 : AOI211_X1 port map( C1 => n2076, C2 => n1373, A => n896, B => n1351,
                           ZN => n899);
   U2529 : INV_X1 port map( A => IRAM_DOUT(5), ZN => n2044);
   U2530 : OAI211_X1 port map( C1 => n1397, C2 => n231, A => n232, B => n233, 
                           ZN => n1537);
   U2531 : NAND4_X1 port map( A1 => n1397, A2 => n1819, A3 => n234, A4 => 
                           IRAM_ADD_9_port, ZN => n232);
   U2532 : AOI21_X1 port map( B1 => n1396, B2 => n1819, A => n236, ZN => n231);
   U2533 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_10_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_10_port, ZN 
                           => n233);
   U2534 : OAI211_X1 port map( C1 => n1395, C2 => n241, A => n242, B => n243, 
                           ZN => n1539);
   U2535 : NAND4_X1 port map( A1 => n1395, A2 => n1819, A3 => n246, A4 => 
                           IRAM_ADD_7_port, ZN => n242);
   U2536 : AOI21_X1 port map( B1 => n1394, B2 => n1819, A => n248, ZN => n241);
   U2537 : AOI22_X1 port map( A1 => n1291, A2 => n191, B1 => n190, B2 => 
                           DATAPATH_IxSecond_stxBR_target_8_port, ZN => n243);
   U2538 : OAI211_X1 port map( C1 => n1393, C2 => n253, A => n254, B => n255, 
                           ZN => n1541);
   U2539 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_6_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_6_port, ZN =>
                           n255);
   U2540 : NAND4_X1 port map( A1 => n1393, A2 => n1819, A3 => n256, A4 => 
                           IRAM_ADD_5_port, ZN => n254);
   U2541 : AOI21_X1 port map( B1 => n1392, B2 => n1819, A => n258, ZN => n253);
   U2542 : OAI211_X1 port map( C1 => n1405, C2 => n187, A => n188, B => n189, 
                           ZN => n1529);
   U2543 : NAND4_X1 port map( A1 => n1405, A2 => n1819, A3 => n192, A4 => 
                           IRAM_ADD_17_port, ZN => n188);
   U2544 : AOI21_X1 port map( B1 => n1404, B2 => n1819, A => n194, ZN => n187);
   U2545 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_18_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_18_port, ZN 
                           => n189);
   U2546 : OAI211_X1 port map( C1 => n1401, C2 => n211, A => n212, B => n213, 
                           ZN => n1533);
   U2547 : NAND4_X1 port map( A1 => n1401, A2 => n1819, A3 => n214, A4 => 
                           IRAM_ADD_13_port, ZN => n212);
   U2548 : AOI21_X1 port map( B1 => n1400, B2 => n1819, A => n216, ZN => n211);
   U2549 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_14_port, B1 => n191, 
                           B2 => DATAPATH_IxSecond_stxjump_target_14_port, ZN 
                           => n213);
   U2550 : OAI211_X1 port map( C1 => n1399, C2 => n221, A => n222, B => n223, 
                           ZN => n1535);
   U2551 : NAND4_X1 port map( A1 => n1399, A2 => n1819, A3 => n224, A4 => 
                           IRAM_ADD_11_port, ZN => n222);
   U2552 : AOI21_X1 port map( B1 => n1398, B2 => n1819, A => n226, ZN => n221);
   U2553 : AOI22_X1 port map( A1 => n190, A2 => 
                           DATAPATH_IxSecond_stxBR_target_12_port, B1 => 
                           DATAPATH_IxSecond_stxjump_target_12_port, B2 => n191
                           , ZN => n223);
   U2554 : NAND2_X1 port map( A1 => n1341, A2 => n1381, ZN => n809);
   U2555 : INV_X1 port map( A => n1047, ZN => n2149);
   U2556 : AOI22_X1 port map( A1 => RF_WR_DATAx15x, A2 => n1577, B1 => 
                           RF_RD2_DATA(15), B2 => n985, ZN => n1048);
   U2557 : INV_X1 port map( A => n1065, ZN => n2156);
   U2558 : OAI21_X1 port map( B1 => n1371, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_15_port);
   U2559 : OAI21_X1 port map( B1 => n1372, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_16_port);
   U2560 : OAI21_X1 port map( B1 => n1373, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_17_port);
   U2561 : OAI21_X1 port map( B1 => n1374, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_18_port);
   U2562 : OAI21_X1 port map( B1 => n1375, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_19_port);
   U2563 : OAI21_X1 port map( B1 => n1376, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_20_port);
   U2564 : OAI21_X1 port map( B1 => n1377, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_21_port);
   U2565 : OAI21_X1 port map( B1 => n1378, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_22_port);
   U2566 : OAI21_X1 port map( B1 => n1379, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_23_port);
   U2567 : OAI21_X1 port map( B1 => n1380, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_24_port);
   U2568 : OAI21_X1 port map( B1 => n1381, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_25_port);
   U2569 : OAI21_X1 port map( B1 => n1382, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_26_port);
   U2570 : OAI21_X1 port map( B1 => n1383, B2 => n1897, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_27_port);
   U2571 : OAI21_X1 port map( B1 => n1384, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_28_port);
   U2572 : OAI21_X1 port map( B1 => n1385, B2 => n963, A => n2092, ZN => 
                           DATAPATH_IxSecond_stximm_extended_30_port);
   U2573 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN2_4_port, ZN => 
                           n1985);
   U2574 : OR2_X1 port map( A1 => n110, A2 => n1416, ZN => n101);
   U2575 : OAI221_X1 port map( B1 => n1860, B2 => n1598, C1 => n1423, C2 => 
                           n1823, A => n1071, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_4_port);
   U2576 : OR3_X1 port map( A1 => n1401, A2 => n1400, A3 => n2205, ZN => n198);
   U2577 : OR3_X1 port map( A1 => n1405, A2 => n1404, A3 => n2204, ZN => n172);
   U2578 : OR3_X1 port map( A1 => n1411, A2 => n1410, A3 => n144, ZN => n132);
   U2579 : OR3_X1 port map( A1 => n1409, A2 => n1408, A3 => n2203, ZN => n144);
   U2580 : INV_X1 port map( A => n945, ZN => n2079);
   U2581 : INV_X1 port map( A => n1028, ZN => RF_WR_DATAx27x);
   U2582 : OAI22_X1 port map( A1 => n1935, A2 => DATAPATH_IxLMD_DATA_27_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_27_port, 
                           ZN => n1028);
   U2583 : INV_X1 port map( A => n1049, ZN => RF_WR_DATAx15x);
   U2584 : OAI22_X1 port map( A1 => n1934, A2 => DATAPATH_IxLMD_DATA_15_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_15_port, 
                           ZN => n1049);
   U2585 : INV_X1 port map( A => n1060, ZN => RF_WR_DATAx11x);
   U2586 : OAI22_X1 port map( A1 => n1933, A2 => DATAPATH_IxLMD_DATA_11_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_11_port, 
                           ZN => n1060);
   U2587 : INV_X1 port map( A => n1039, ZN => RF_WR_DATAx8x);
   U2588 : OAI22_X1 port map( A1 => n1935, A2 => DATAPATH_IxLMD_DATA_8_port, B1
                           => n1931, B2 => DATAPATH_IxALUOUT_Data1_8_port, ZN 
                           => n1039);
   U2589 : INV_X1 port map( A => n1025, ZN => RF_WR_DATAx26x);
   U2590 : OAI22_X1 port map( A1 => n1935, A2 => DATAPATH_IxLMD_DATA_26_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_26_port, 
                           ZN => n1025);
   U2591 : INV_X1 port map( A => n1045, ZN => RF_WR_DATAx14x);
   U2592 : OAI22_X1 port map( A1 => n1934, A2 => DATAPATH_IxLMD_DATA_14_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_14_port, 
                           ZN => n1045);
   U2593 : INV_X1 port map( A => n1053, ZN => RF_WR_DATAx12x);
   U2594 : OAI22_X1 port map( A1 => n1934, A2 => DATAPATH_IxLMD_DATA_12_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_12_port, 
                           ZN => n1053);
   U2595 : INV_X1 port map( A => n1042, ZN => RF_WR_DATAx9x);
   U2596 : OAI22_X1 port map( A1 => n1934, A2 => DATAPATH_IxLMD_DATA_9_port, B1
                           => n1931, B2 => DATAPATH_IxALUOUT_Data1_9_port, ZN 
                           => n1042);
   U2597 : INV_X1 port map( A => n1034, ZN => RF_WR_DATAx29x);
   U2598 : OAI22_X1 port map( A1 => n1935, A2 => DATAPATH_IxLMD_DATA_29_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_29_port, 
                           ZN => n1034);
   U2599 : INV_X1 port map( A => n1082, ZN => RF_WR_DATAx2x);
   U2600 : OAI22_X1 port map( A1 => n1932, A2 => DATAPATH_IxLMD_DATA_2_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_2_port, ZN 
                           => n1082);
   U2601 : INV_X1 port map( A => n1070, ZN => RF_WR_DATAx0x);
   U2602 : OAI22_X1 port map( A1 => n1933, A2 => DATAPATH_IxLMD_DATA_0_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_0_port, ZN 
                           => n1070);
   U2603 : INV_X1 port map( A => n1085, ZN => RF_WR_DATAx3x);
   U2604 : OAI22_X1 port map( A1 => n1932, A2 => DATAPATH_IxLMD_DATA_3_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_3_port, ZN 
                           => n1085);
   U2605 : INV_X1 port map( A => n1114, ZN => RF_WR_DATAx1x);
   U2606 : OAI22_X1 port map( A1 => n1932, A2 => DATAPATH_IxLMD_DATA_1_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_1_port, ZN 
                           => n1114);
   U2607 : INV_X1 port map( A => n1067, ZN => RF_WR_DATAx7x);
   U2608 : OAI22_X1 port map( A1 => n1933, A2 => DATAPATH_IxLMD_DATA_7_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_7_port, ZN 
                           => n1067);
   U2609 : INV_X1 port map( A => n1079, ZN => RF_WR_DATAx6x);
   U2610 : OAI22_X1 port map( A1 => n1932, A2 => DATAPATH_IxLMD_DATA_6_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_6_port, ZN 
                           => n1079);
   U2611 : INV_X1 port map( A => n1073, ZN => RF_WR_DATAx4x);
   U2612 : OAI22_X1 port map( A1 => n1933, A2 => DATAPATH_IxLMD_DATA_4_port, B1
                           => n1590, B2 => DATAPATH_IxALUOUT_Data1_4_port, ZN 
                           => n1073);
   U2613 : INV_X1 port map( A => n1018, ZN => RF_WR_DATAx25x);
   U2614 : OAI22_X1 port map( A1 => n1936, A2 => DATAPATH_IxLMD_DATA_25_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_25_port, 
                           ZN => n1018);
   U2615 : INV_X1 port map( A => n986, ZN => RF_WR_DATAx19x);
   U2616 : OAI22_X1 port map( A1 => n1938, A2 => DATAPATH_IxLMD_DATA_19_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_19_port, 
                           ZN => n986);
   U2617 : INV_X1 port map( A => n1003, ZN => RF_WR_DATAx23x);
   U2618 : OAI22_X1 port map( A1 => n1937, A2 => DATAPATH_IxLMD_DATA_23_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_23_port, 
                           ZN => n1003);
   U2619 : INV_X1 port map( A => n996, ZN => RF_WR_DATAx20x);
   U2620 : OAI22_X1 port map( A1 => n1937, A2 => DATAPATH_IxLMD_DATA_20_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_20_port, 
                           ZN => n996);
   U2621 : INV_X1 port map( A => n1015, ZN => RF_WR_DATAx31x);
   U2622 : OAI22_X1 port map( A1 => n1936, A2 => DATAPATH_IxLMD_DATA_31_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_31_port, 
                           ZN => n1015);
   U2623 : INV_X1 port map( A => n993, ZN => RF_WR_DATAx16x);
   U2624 : OAI22_X1 port map( A1 => n1937, A2 => DATAPATH_IxLMD_DATA_16_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_16_port, 
                           ZN => n993);
   U2625 : INV_X1 port map( A => n1009, ZN => RF_WR_DATAx17x);
   U2626 : OAI22_X1 port map( A1 => n1936, A2 => DATAPATH_IxLMD_DATA_17_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_17_port, 
                           ZN => n1009);
   U2627 : INV_X1 port map( A => n1006, ZN => RF_WR_DATAx18x);
   U2628 : OAI22_X1 port map( A1 => n1937, A2 => DATAPATH_IxLMD_DATA_18_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_18_port, 
                           ZN => n1006);
   U2629 : INV_X1 port map( A => n999, ZN => RF_WR_DATAx21x);
   U2630 : OAI22_X1 port map( A1 => n1937, A2 => DATAPATH_IxLMD_DATA_21_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_21_port, 
                           ZN => n999);
   U2631 : INV_X1 port map( A => n990, ZN => RF_WR_DATAx22x);
   U2632 : OAI22_X1 port map( A1 => n1938, A2 => DATAPATH_IxLMD_DATA_22_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_22_port, 
                           ZN => n990);
   U2633 : INV_X1 port map( A => n1063, ZN => RF_WR_DATAx13x);
   U2634 : OAI22_X1 port map( A1 => n1933, A2 => DATAPATH_IxLMD_DATA_13_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_13_port, 
                           ZN => n1063);
   U2635 : INV_X1 port map( A => n1056, ZN => RF_WR_DATAx10x);
   U2636 : OAI22_X1 port map( A1 => n1934, A2 => DATAPATH_IxLMD_DATA_10_port, 
                           B1 => n1931, B2 => DATAPATH_IxALUOUT_Data1_10_port, 
                           ZN => n1056);
   U2637 : INV_X1 port map( A => n1012, ZN => RF_WR_DATAx30x);
   U2638 : OAI22_X1 port map( A1 => n1936, A2 => DATAPATH_IxLMD_DATA_30_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_30_port, 
                           ZN => n1012);
   U2639 : INV_X1 port map( A => n1021, ZN => RF_WR_DATAx24x);
   U2640 : OAI22_X1 port map( A1 => n1936, A2 => DATAPATH_IxLMD_DATA_24_port, 
                           B1 => n1590, B2 => DATAPATH_IxALUOUT_Data1_24_port, 
                           ZN => n1021);
   U2641 : OAI221_X1 port map( B1 => n1861, B2 => n1616, C1 => n1449, C2 => 
                           n1950, A => n1010, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_30_port);
   U2642 : INV_X1 port map( A => IRAM_DOUT(1), ZN => n2047);
   U2643 : INV_X1 port map( A => IRAM_DOUT(0), ZN => n2048);
   U2644 : OR3_X1 port map( A1 => IRAM_DOUT(2), A2 => IRAM_DOUT(5), A3 => n2042
                           , ZN => n1139);
   U2645 : OAI221_X1 port map( B1 => n1880, B2 => n1617, C1 => n1442, C2 => 
                           n1950, A => n1000, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_23_port);
   U2646 : AND2_X1 port map( A1 => CU_Ixcw2_i_11_port, A2 => n1750, ZN => n1864
                           );
   U2647 : NOR3_X1 port map( A1 => n1336, A2 => n1335, A3 => n1918, ZN => n334)
                           ;
   U2648 : XNOR2_X1 port map( A => n1361, B => n1386, ZN => n839);
   U2649 : XNOR2_X1 port map( A => n1357, B => n1386, ZN => n855);
   U2650 : XNOR2_X1 port map( A => n1356, B => n1386, ZN => n854);
   U2651 : XNOR2_X1 port map( A => n1360, B => n1386, ZN => n838);
   U2652 : NOR2_X1 port map( A1 => n1385, A2 => n1345, ZN => n933);
   U2653 : NOR3_X1 port map( A1 => n2004, A2 => IRAM_DOUT(14), A3 => 
                           IRAM_DOUT(12), ZN => n38);
   U2654 : AOI21_X1 port map( B1 => n1362, B2 => n1363, A => n1386, ZN => n824)
                           ;
   U2655 : AOI21_X1 port map( B1 => n1358, B2 => n1359, A => n1386, ZN => n843)
                           ;
   U2656 : AOI21_X1 port map( B1 => n1354, B2 => n1355, A => n1386, ZN => n860)
                           ;
   U2657 : XNOR2_X1 port map( A => n1355, B => n1914, ZN => n852);
   U2658 : XNOR2_X1 port map( A => n1359, B => n1914, ZN => n836);
   U2659 : OAI22_X1 port map( A1 => n1276, A2 => n1993, B1 => n1335, B2 => 
                           n1991, ZN => n1286);
   U2660 : OAI22_X1 port map( A1 => n1275, A2 => n1993, B1 => n1336, B2 => 
                           n1991, ZN => n1285);
   U2661 : OAI22_X1 port map( A1 => n1298, A2 => n1706, B1 => n1133, B2 => n26,
                           ZN => CU_IxN51);
   U2662 : OAI22_X1 port map( A1 => n1298, A2 => n1706, B1 => n1133, B2 => 
                           n1134, ZN => CU_IxN52);
   U2663 : OAI21_X1 port map( B1 => n1359, B2 => n1358, A => n1386, ZN => n845)
                           ;
   U2664 : OAI21_X1 port map( B1 => n1355, B2 => n1354, A => n1386, ZN => n862)
                           ;
   U2665 : OAI21_X1 port map( B1 => n1363, B2 => n1362, A => n1386, ZN => n826)
                           ;
   U2666 : OAI22_X1 port map( A1 => n1274, A2 => n1993, B1 => n1921, B2 => 
                           n1991, ZN => n1284);
   U2667 : NOR2_X1 port map( A1 => n1197, A2 => n298, ZN => n1133);
   U2668 : XNOR2_X1 port map( A => n1358, B => n1915, ZN => n152);
   U2669 : XNOR2_X1 port map( A => n1354, B => n1915, ZN => n180);
   U2670 : NOR3_X1 port map( A1 => n2004, A2 => IRAM_DOUT(5), A3 => 
                           IRAM_DOUT(2), ZN => n43);
   U2671 : XNOR2_X1 port map( A => n2033, B => IRAM_DOUT(13), ZN => n29);
   U2672 : OR2_X1 port map( A1 => n1929, A2 => n1336, ZN => n1865);
   U2673 : NAND2_X1 port map( A1 => n1344, A2 => n1646, ZN => n950);
   U2674 : AND2_X1 port map( A1 => n1345, A2 => n1385, ZN => n941);
   U2675 : NAND2_X1 port map( A1 => n950, A2 => n951, ZN => n946);
   U2676 : AND2_X1 port map( A1 => n1382, A2 => n1342, ZN => n801);
   U2677 : INV_X1 port map( A => IRAM_DOUT(14), ZN => n2033);
   U2678 : INV_X1 port map( A => n35, ZN => n2003);
   U2679 : OAI22_X1 port map( A1 => n26, A2 => n1993, B1 => n1991, B2 => n1275,
                           ZN => n35);
   U2680 : INV_X1 port map( A => IRAM_DOUT(12), ZN => n2035);
   U2681 : AOI22_X1 port map( A1 => n37, A2 => n38, B1 => n1993, B2 => n1642, 
                           ZN => n36);
   U2682 : NOR2_X1 port map( A1 => n2044, A2 => n2034, ZN => n37);
   U2683 : INV_X1 port map( A => n25, ZN => n2002);
   U2684 : NAND4_X1 port map( A1 => n27, A2 => n28, A3 => n29, A4 => n2035, ZN 
                           => n22);
   U2685 : OAI22_X1 port map( A1 => n26, A2 => n1993, B1 => n1991, B2 => n1274,
                           ZN => n25);
   U2686 : INV_X1 port map( A => IRAM_DOUT(13), ZN => n2034);
   U2687 : OR2_X1 port map( A1 => n32, A2 => IRAM_DOUT(13), ZN => n23);
   U2688 : INV_X1 port map( A => n1881, ZN => n1866);
   U2689 : INV_X1 port map( A => n1587, ZN => n2106);
   U2690 : AOI21_X1 port map( B1 => n1957, B2 => n1784, A => n1955, ZN => n516)
                           ;
   U2691 : NOR2_X1 port map( A1 => n1785, A2 => n495, ZN => n497);
   U2692 : AOI22_X1 port map( A1 => RF_WR_DATAx6x, A2 => n1578, B1 => 
                           RF_RD2_DATA(6), B2 => n1940, ZN => n1078);
   U2693 : AOI22_X1 port map( A1 => RF_WR_DATAx5x, A2 => n1578, B1 => 
                           RF_RD2_DATA(5), B2 => n1816, ZN => n1075);
   U2694 : AOI22_X1 port map( A1 => RF_WR_DATAx4x, A2 => n1578, B1 => 
                           RF_RD2_DATA(4), B2 => n1816, ZN => n1072);
   U2695 : AOI22_X1 port map( A1 => RF_WR_DATAx7x, A2 => n1578, B1 => 
                           RF_RD2_DATA(7), B2 => n985, ZN => n1066);
   U2696 : AOI22_X1 port map( A1 => n1578, A2 => RF_WR_DATAx2x, B1 => 
                           RF_RD2_DATA(2), B2 => n985, ZN => n1081);
   U2697 : AOI22_X1 port map( A1 => RF_WR_DATAx1x, A2 => n1943, B1 => 
                           RF_RD2_DATA(1), B2 => n1940, ZN => n1109);
   U2698 : AOI21_X1 port map( B1 => n767, B2 => n689, A => n677, ZN => n766);
   U2699 : XNOR2_X1 port map( A => n2117, B => n664, ZN => n661);
   U2700 : AOI21_X1 port map( B1 => n647, B2 => n2117, A => n649, ZN => n656);
   U2701 : INV_X1 port map( A => n1759, ZN => n2089);
   U2702 : OAI21_X1 port map( B1 => n270, B2 => n1729, A => n2084, ZN => n812);
   U2703 : OAI21_X1 port map( B1 => n1386, B2 => n2057, A => n1358, ZN => n849)
                           ;
   U2704 : AOI21_X1 port map( B1 => n696, B2 => n1928, A => n1652, ZN => n781);
   U2705 : OAI211_X1 port map( C1 => n1768, C2 => n2161, A => n699, B => n698, 
                           ZN => DATAPATH_IxThird_stxALU_out_i_0_port);
   U2706 : AOI22_X1 port map( A1 => n703, A2 => n702, B1 => n2129, B2 => n1990,
                           ZN => n698);
   U2707 : XNOR2_X1 port map( A => n1920, B => 
                           DATAPATH_IxThird_stxALU_IN2_0_port, ZN => n569);
   U2708 : INV_X1 port map( A => n111, ZN => n2061);
   U2709 : AOI21_X1 port map( B1 => n718, B2 => n433, A => n719, ZN => n716);
   U2710 : OAI221_X1 port map( B1 => n1235, B2 => n1906, C1 => n111, C2 => 
                           n1904, A => n112, ZN => n1518);
   U2711 : XNOR2_X1 port map( A => n831, B => n830, ZN => n111);
   U2712 : AOI21_X1 port map( B1 => RF_RD1_ADD_4_port, B2 => n1764, A => n882, 
                           ZN => n867);
   U2713 : NOR2_X1 port map( A1 => n1764, A2 => n882, ZN => n896);
   U2714 : NOR2_X1 port map( A1 => n1764, A2 => n1386, ZN => n882);
   U2715 : AOI21_X1 port map( B1 => n759, B2 => n645, A => n633, ZN => n758);
   U2716 : NAND2_X1 port map( A1 => n1780, A2 => CU_Ixcw2_i_12_port, ZN => n897
                           );
   U2717 : AOI21_X1 port map( B1 => n780, B2 => n1710, A => n407, ZN => n779);
   U2718 : AND2_X1 port map( A1 => CU_Ixcw_LUT_0_port, A2 => n1842, ZN => 
                           CU_Ixcw1_0_port);
   U2719 : AND2_X1 port map( A1 => CU_Ixcw_LUT_10_port, A2 => n1842, ZN => 
                           CU_Ixcw1_10_port);
   U2720 : AND2_X1 port map( A1 => CU_Ixcw_LUT_1_port, A2 => n1842, ZN => 
                           CU_Ixcw1_1_port);
   U2721 : AND2_X1 port map( A1 => CU_Ixcw_LUT_2_port, A2 => n1842, ZN => 
                           CU_Ixcw1_2_port);
   U2722 : AND2_X1 port map( A1 => CU_Ixcw_LUT_4_port, A2 => n1842, ZN => 
                           CU_Ixcw1_4_port);
   U2723 : AND2_X1 port map( A1 => CU_Ixcw_LUT_5_port, A2 => n1842, ZN => 
                           CU_Ixcw1_5_port);
   U2724 : AND2_X1 port map( A1 => CU_Ixcw_LUT_7_port, A2 => n1842, ZN => 
                           CU_Ixcw1_7_port);
   U2725 : AND2_X1 port map( A1 => CU_Ixcw_LUT_8_port, A2 => n1842, ZN => 
                           CU_Ixcw1_8_port);
   U2726 : AND2_X1 port map( A1 => CU_Ixcw_LUT_6_port, A2 => n1842, ZN => 
                           CU_Ixcw1_6_port);
   U2727 : AND2_X1 port map( A1 => CU_Ixcw_LUT_9_port, A2 => n1842, ZN => 
                           CU_Ixcw1_9_port);
   U2728 : AOI21_X1 port map( B1 => n739, B2 => n491, A => n478, ZN => n738);
   U2729 : NAND2_X1 port map( A1 => n1849, A2 => n1991, ZN => n92);
   U2730 : NOR2_X1 port map( A1 => CU_Ixcw_LUT_16_port, A2 => n1849, ZN => 
                           CU_Ixcw1_14_port);
   U2731 : AOI21_X1 port map( B1 => n746, B2 => n539, A => n527, ZN => n745);
   U2732 : CLKBUF_X1 port map( A => n1751, Z => n1867);
   U2733 : OAI22_X1 port map( A1 => n2122, A2 => n773, B1 => n774, B2 => n359, 
                           ZN => n338);
   U2734 : AOI22_X1 port map( A1 => n1909, A2 => n565, B1 => 
                           DATAPATH_IxThird_stxALU1xN192, B2 => n1958, ZN => 
                           n564);
   U2735 : INV_X1 port map( A => n1838, ZN => n2114);
   U2736 : NAND2_X1 port map( A1 => n601, A2 => n1838, ZN => n613);
   U2737 : AOI22_X1 port map( A1 => n2114, A2 => n595, B1 => n596, B2 => n1838,
                           ZN => n590);
   U2738 : AOI22_X1 port map( A1 => n2114, A2 => n578, B1 => n579, B2 => n1838,
                           ZN => n572);
   U2739 : XNOR2_X1 port map( A => n1922, B => n1679, ZN => n582);
   U2740 : AOI22_X1 port map( A1 => n1909, A2 => n1679, B1 => 
                           DATAPATH_IxThird_stxALU1xN210, B2 => n1958, ZN => 
                           n575);
   U2741 : INV_X1 port map( A => n283, ZN => n2091);
   U2742 : OR2_X2 port map( A1 => n1088, A2 => n1090, ZN => n1876);
   U2743 : INV_X1 port map( A => n1881, ZN => n981);
   U2744 : BUF_X2 port map( A => n1891, Z => n1947);
   U2745 : OR2_X2 port map( A1 => n1088, A2 => n2201, ZN => n1879);
   U2746 : BUF_X1 port map( A => n1876, Z => n1880);
   U2747 : INV_X2 port map( A => n1879, ZN => n1948);
   U2748 : NAND2_X1 port map( A1 => n1094, A2 => n1095, ZN => n1092);
   U2749 : INV_X1 port map( A => n1113, ZN => n2200);
   U2750 : OAI221_X1 port map( B1 => n1911, B2 => n514, C1 => n2140, C2 => n516
                           , A => n517, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_23_port);
   U2751 : XNOR2_X1 port map( A => n1918, B => n2140, ZN => n744);
   U2752 : INV_X1 port map( A => n1001, ZN => n2140);
   U2753 : INV_X1 port map( A => n1734, ZN => n2127);
   U2754 : NOR4_X1 port map( A1 => n565, A2 => n399, A3 => n790, A4 => n1656, 
                           ZN => n967);
   U2755 : AND2_X1 port map( A1 => n1113, A2 => n1111, ZN => n1881);
   U2756 : NOR4_X1 port map( A1 => n1893, A2 => n1894, A3 => n1895, A4 => n1896
                           , ZN => n1882);
   U2757 : XNOR2_X1 port map( A => n1883, B => n1159, ZN => n1131);
   U2758 : AND3_X1 port map( A1 => n1952, A2 => n1879, A3 => n1876, ZN => n1884
                           );
   U2759 : CLKBUF_X1 port map( A => n536, Z => n1885);
   U2760 : CLKBUF_X1 port map( A => n1671, Z => n1886);
   U2761 : NOR2_X1 port map( A1 => n487, A2 => n469, ZN => n1022);
   U2762 : XNOR2_X1 port map( A => n1918, B => n1805, ZN => n491);
   U2763 : NOR4_X1 port map( A1 => n1097, A2 => n1334, A3 => n1882, A4 => n1333
                           , ZN => n1095);
   U2764 : NOR4_X1 port map( A1 => n1893, A2 => n1894, A3 => n1896, A4 => n1895
                           , ZN => n1096);
   U2765 : XNOR2_X1 port map( A => n1887, B => n1160, ZN => n1130);
   U2766 : XNOR2_X1 port map( A => n2151, B => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, ZN => n655);
   U2767 : OAI221_X1 port map( B1 => n1432, B2 => n1762, C1 => n1188, C2 => 
                           n1769, A => n1062, ZN => n762);
   U2768 : AOI22_X1 port map( A1 => RF_WR_DATAx13x, A2 => n1578, B1 => 
                           RF_RD2_DATA(13), B2 => n985, ZN => n1062);
   U2769 : AOI22_X1 port map( A1 => n1910, A2 => n1801, B1 => 
                           DATAPATH_IxThird_stxALU1xN201, B2 => n1958, ZN => 
                           n685);
   U2770 : XNOR2_X1 port map( A => n1919, B => n1801, ZN => n689);
   U2771 : AND3_X1 port map( A1 => n1952, A2 => n1879, A3 => n1876, ZN => n1888
                           );
   U2772 : OAI221_X1 port map( B1 => n2130, B2 => n416, C1 => n2049, C2 => n418
                           , A => n419, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_31_port);
   U2773 : XNOR2_X1 port map( A => n2130, B => DATAPATH_IxThird_stxALU1xN222, 
                           ZN => n422);
   U2774 : INV_X1 port map( A => n715, ZN => n2130);
   U2775 : OAI221_X1 port map( B1 => n1434, B2 => n1762, C1 => n1181, C2 => 
                           n1869, A => n1048, ZN => n1047);
   U2776 : AOI22_X1 port map( A1 => n1909, A2 => n610, B1 => 
                           DATAPATH_IxThird_stxALU1xN208, B2 => n1959, ZN => 
                           n609);
   U2777 : XNOR2_X1 port map( A => n2146, B => 
                           DATAPATH_IxThird_stxALU_IN1_17_port, ZN => n610);
   U2778 : INV_X1 port map( A => n787, ZN => n2146);
   U2779 : XNOR2_X1 port map( A => n1919, B => n1582, ZN => n605);
   U2780 : OAI221_X1 port map( B1 => n1436, B2 => n1761, C1 => n1176, C2 => 
                           n1869, A => n1008, ZN => n787);
   U2781 : XNOR2_X1 port map( A => n2138, B => 
                           DATAPATH_IxThird_stxALU_IN1_24_port, ZN => n512);
   U2782 : XNOR2_X1 port map( A => n1920, B => n762, ZN => n650);
   U2783 : INV_X1 port map( A => n762, ZN => n2151);
   U2784 : OAI221_X1 port map( B1 => n2142, B2 => n548, C1 => n1912, C2 => n549
                           , A => n550, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_21_port);
   U2785 : AOI22_X1 port map( A1 => n1909, A2 => n1588, B1 => 
                           DATAPATH_IxThird_stxALU1xN211, B2 => n1959, ZN => 
                           n559);
   U2786 : XNOR2_X1 port map( A => n1918, B => n1588, ZN => n561);
   U2787 : XNOR2_X1 port map( A => n1920, B => n750, ZN => n543);
   U2788 : INV_X1 port map( A => n750, ZN => n2143);
   U2789 : AOI22_X1 port map( A1 => n1909, A2 => n1672, B1 => 
                           DATAPATH_IxThird_stxALU1xN209, B2 => n1958, ZN => 
                           n593);
   U2790 : OAI221_X1 port map( B1 => n1437, B2 => n1762, C1 => n1175, C2 => 
                           n1868, A => n1005, ZN => n785);
   U2791 : XNOR2_X1 port map( A => n2141, B => 
                           DATAPATH_IxThird_stxALU_IN1_22_port, ZN => n536);
   U2792 : OAI221_X1 port map( B1 => n1911, B2 => n532, C1 => n2141, C2 => n534
                           , A => n535, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_22_port);
   U2793 : INV_X1 port map( A => n980, ZN => n1889);
   U2794 : BUF_X2 port map( A => n1808, Z => n1940);
   U2795 : OAI221_X1 port map( B1 => n2147, B2 => n615, C1 => n1913, C2 => n616
                           , A => n617, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_16_port);
   U2796 : XNOR2_X1 port map( A => n1918, B => n788, ZN => n601);
   U2797 : XNOR2_X1 port map( A => n2137, B => 
                           DATAPATH_IxThird_stxALU_IN1_25_port, ZN => n503);
   U2798 : INV_X1 port map( A => n741, ZN => n2137);
   U2799 : OAI221_X1 port map( B1 => n1444, B2 => n1761, C1 => n1171, C2 => 
                           n1769, A => n1017, ZN => n741);
   U2800 : AOI22_X1 port map( A1 => n1910, A2 => n1725, B1 => 
                           DATAPATH_IxThird_stxALU1xN202, B2 => n1958, ZN => 
                           n668);
   U2801 : XNOR2_X1 port map( A => n1927, B => n1725, ZN => n674);
   U2802 : XNOR2_X1 port map( A => n1918, B => n749, ZN => n546);
   U2803 : XNOR2_X1 port map( A => n1923, B => n1988, ZN => n413);
   U2804 : AND4_X1 port map( A1 => n1155, A2 => n1156, A3 => n1154, A4 => n1132
                           , ZN => n1120);
   U2805 : AOI22_X1 port map( A1 => n1910, A2 => n642, B1 => 
                           DATAPATH_IxThird_stxALU1xN205, B2 => n1958, ZN => 
                           n641);
   U2806 : XNOR2_X1 port map( A => n1919, B => n642, ZN => n645);
   U2807 : XNOR2_X1 port map( A => n2150, B => 
                           DATAPATH_IxThird_stxALU_IN1_14_port, ZN => n642);
   U2808 : XNOR2_X1 port map( A => n1927, B => n760, ZN => n636);
   U2809 : AOI22_X1 port map( A1 => n1908, A2 => n1802, B1 => 
                           DATAPATH_IxThird_stxALU1xN221, B2 => n1959, ZN => 
                           n426);
   U2810 : XNOR2_X1 port map( A => n1918, B => n1802, ZN => n433);
   U2811 : XNOR2_X1 port map( A => n1918, B => n731, ZN => n730);
   U2812 : AOI22_X1 port map( A1 => n1909, A2 => n1721, B1 => 
                           DATAPATH_IxThird_stxALU1xN207, B2 => n1958, ZN => 
                           n617);
   U2813 : XNOR2_X1 port map( A => n1926, B => n1721, ZN => n619);
   U2814 : XNOR2_X1 port map( A => n1919, B => n1889, ZN => n753);
   U2815 : NAND2_X1 port map( A1 => n1118, A2 => n1119, ZN => n1116);
   U2816 : AND3_X1 port map( A1 => n1952, A2 => n1879, A3 => n1876, ZN => n1890
                           );
   U2817 : CLKBUF_X1 port map( A => n1884, Z => n1946);
   U2818 : CLKBUF_X1 port map( A => n2077, Z => n1892);
   U2819 : OAI21_X1 port map( B1 => n1754, B2 => IMM_SEL_i, A => n1116, ZN => 
                           n1111);
   U2820 : XNOR2_X1 port map( A => n2153, B => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, ZN => n686);
   U2821 : INV_X1 port map( A => n768, ZN => n2153);
   U2822 : AOI22_X1 port map( A1 => RF_WR_DATAx10x, A2 => n1578, B1 => 
                           RF_RD2_DATA(10), B2 => n985, ZN => n1055);
   U2823 : XNOR2_X1 port map( A => n1158, B => n1154, ZN => n1126);
   U2824 : XNOR2_X1 port map( A => n2145, B => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, ZN => n594);
   U2825 : INV_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_18_port, ZN => 
                           n2111);
   U2826 : XNOR2_X1 port map( A => n1918, B => n1672, ZN => n597);
   U2827 : XNOR2_X1 port map( A => n1922, B => n785, ZN => n588);
   U2828 : OAI221_X1 port map( B1 => n1425, B2 => n1761, C1 => n1190, C2 => 
                           n1869, A => n1078, ZN => n372);
   U2829 : OAI221_X1 port map( B1 => n1424, B2 => n1762, C1 => n1191, C2 => 
                           n1770, A => n1075, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_5_port);
   U2830 : OAI221_X1 port map( B1 => n1423, B2 => n1762, C1 => n1192, C2 => 
                           n1769, A => n1072, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_4_port);
   U2831 : OAI221_X1 port map( B1 => n1420, B2 => n1761, C1 => n1194, C2 => 
                           n1769, A => n1109, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_1_port);
   U2832 : OAI221_X1 port map( B1 => n1426, B2 => n1762, C1 => n1189, C2 => 
                           n1770, A => n1066, ZN => n1065);
   U2833 : OAI221_X1 port map( B1 => n1421, B2 => n1762, C1 => n1195, C2 => 
                           n1868, A => n1081, ZN => 
                           DATAPATH_IxThird_stxALU_IN2_2_port);
   U2834 : INV_X1 port map( A => n1843, ZN => n2099);
   U2835 : XNOR2_X1 port map( A => n1918, B => n1843, ZN => n464);
   U2836 : NAND2_X1 port map( A1 => n1877, A2 => n1878, ZN => n1896);
   U2837 : XNOR2_X1 port map( A => n2131, B => 
                           DATAPATH_IxThird_stxALU_IN1_30_port, ZN => n427);
   U2838 : INV_X1 port map( A => n731, ZN => n2131);
   U2839 : AOI22_X1 port map( A1 => RF_WR_DATAx24x, A2 => n1943, B1 => 
                           RF_RD2_DATA(24), B2 => n1941, ZN => n1020);
   U2840 : AOI22_X1 port map( A1 => RF_WR_DATAx17x, A2 => n1578, B1 => 
                           RF_RD2_DATA(17), B2 => n1941, ZN => n1008);
   U2841 : AOI22_X1 port map( A1 => RF_WR_DATAx20x, A2 => n1578, B1 => 
                           RF_RD2_DATA(20), B2 => n1940, ZN => n995);
   U2842 : AOI22_X1 port map( A1 => RF_WR_DATAx25x, A2 => n1943, B1 => 
                           RF_RD2_DATA(25), B2 => n985, ZN => n1017);
   U2843 : AOI22_X1 port map( A1 => RF_WR_DATAx31x, A2 => n1943, B1 => 
                           RF_RD2_DATA(31), B2 => n1816, ZN => n1014);
   U2844 : AOI22_X1 port map( A1 => RF_WR_DATAx16x, A2 => n1943, B1 => 
                           RF_RD2_DATA(16), B2 => n1940, ZN => n992);
   U2845 : AOI22_X1 port map( A1 => RF_WR_DATAx18x, A2 => n1578, B1 => 
                           RF_RD2_DATA(18), B2 => n1940, ZN => n1005);
   U2846 : AOI22_X1 port map( A1 => RF_WR_DATAx30x, A2 => n1943, B1 => 
                           RF_RD2_DATA(30), B2 => n1816, ZN => n1011);
   U2847 : AOI22_X1 port map( A1 => RF_WR_DATAx22x, A2 => n1943, B1 => 
                           RF_RD2_DATA(22), B2 => n1816, ZN => n989);
   U2848 : XNOR2_X1 port map( A => n1153, B => n1146, ZN => n1128);
   U2849 : XNOR2_X1 port map( A => n1795, B => 
                           DATAPATH_IxThird_stxALU_IN1_23_port, ZN => n518);
   U2850 : OAI221_X1 port map( B1 => n1442, B2 => n1762, C1 => n1174, C2 => 
                           n1868, A => n1002, ZN => n1001);
   U2851 : AOI22_X1 port map( A1 => RF_WR_DATAx23x, A2 => n1578, B1 => 
                           RF_RD2_DATA(23), B2 => n1816, ZN => n1002);
   U2852 : AOI22_X1 port map( A1 => RF_WR_DATAx5x, A2 => n1948, B1 => 
                           RF_RD1_DATA(5), B2 => n1946, ZN => n1074);
   U2853 : AOI22_X1 port map( A1 => RF_WR_DATAx3x, A2 => n1948, B1 => 
                           RF_RD1_DATA(3), B2 => n1947, ZN => n1083);
   U2854 : AOI22_X1 port map( A1 => RF_WR_DATAx4x, A2 => n1948, B1 => 
                           RF_RD1_DATA(4), B2 => n1946, ZN => n1071);
   U2855 : AOI22_X1 port map( A1 => RF_WR_DATAx6x, A2 => n1948, B1 => 
                           RF_RD1_DATA(6), B2 => n1947, ZN => n1077);
   U2856 : AOI22_X1 port map( A1 => RF_WR_DATAx0x, A2 => n1948, B1 => 
                           RF_RD1_DATA(0), B2 => n1947, ZN => n1068);
   U2857 : AOI22_X1 port map( A1 => n1948, A2 => RF_WR_DATAx2x, B1 => 
                           RF_RD1_DATA(2), B2 => n1947, ZN => n1080);
   U2858 : AOI22_X1 port map( A1 => RF_WR_DATAx7x, A2 => n1948, B1 => 
                           RF_RD1_DATA(7), B2 => n1888, ZN => n1064);
   U2859 : AOI22_X1 port map( A1 => RF_RD1_DATA(29), A2 => n1890, B1 => 
                           RF_WR_DATAx29x, B2 => n1948, ZN => n1032);
   U2860 : AOI22_X1 port map( A1 => RF_WR_DATAx12x, A2 => n1948, B1 => 
                           RF_RD1_DATA(12), B2 => n979, ZN => n1050);
   U2861 : AOI22_X1 port map( A1 => RF_WR_DATAx10x, A2 => n1948, B1 => 
                           RF_RD1_DATA(10), B2 => n1890, ZN => n1054);
   U2862 : NOR4_X1 port map( A1 => n1106, A2 => n1096, A3 => n1107, A4 => n1299
                           , ZN => n1105);
   U2863 : INV_X1 port map( A => n749, ZN => n2142);
   U2864 : AOI22_X1 port map( A1 => RF_WR_DATAx21x, A2 => n1578, B1 => 
                           RF_RD2_DATA(21), B2 => n1940, ZN => n998);
   U2865 : OAI221_X4 port map( B1 => n1871, B2 => n1612, C1 => n1439, C2 => 
                           n1950, A => n994, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_20_port);
   U2866 : AOI21_X1 port map( B1 => n1755, B2 => n2084, A => n270, ZN => n954);
   U2867 : AOI22_X1 port map( A1 => n1909, A2 => n1650, B1 => 
                           DATAPATH_IxThird_stxALU1xN214, B2 => n1959, ZN => 
                           n517);
   U2868 : XNOR2_X1 port map( A => n1925, B => n518, ZN => n524);
   U2869 : XNOR2_X1 port map( A => n1152, B => n1145, ZN => n1127);
   U2870 : AND2_X1 port map( A1 => n1152, A2 => n1153, ZN => n1132);
   U2871 : AOI21_X1 port map( B1 => n1956, B2 => n1663, A => n1955, ZN => n574)
                           ;
   U2872 : INV_X1 port map( A => n1663, ZN => n2110);
   U2873 : OAI221_X1 port map( B1 => n1880, B2 => n1600, C1 => n1438, C2 => 
                           n1950, A => n977, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_19_port);
   U2874 : AOI22_X1 port map( A1 => RF_WR_DATAx19x, A2 => n1948, B1 => n1884, 
                           B2 => RF_RD1_DATA(19), ZN => n977);
   U2875 : AOI22_X1 port map( A1 => n1909, A2 => n1885, B1 => 
                           DATAPATH_IxThird_stxALU1xN213, B2 => n1959, ZN => 
                           n535);
   U2876 : XNOR2_X1 port map( A => n1918, B => n1885, ZN => n539);
   U2877 : XNOR2_X1 port map( A => n1926, B => n747, ZN => n530);
   U2878 : INV_X1 port map( A => n747, ZN => n2141);
   U2879 : NAND2_X1 port map( A1 => n1115, A2 => n1116, ZN => n1113);
   U2880 : AOI21_X1 port map( B1 => n953, B2 => n808, A => n805, ZN => n952);
   U2881 : OAI21_X1 port map( B1 => n954, B2 => n813, A => n2199, ZN => n953);
   U2882 : OAI221_X1 port map( B1 => n1438, B2 => n1761, C1 => n1177, C2 => 
                           n1869, A => n983, ZN => n980);
   U2883 : AOI22_X1 port map( A1 => RF_WR_DATAx19x, A2 => n1578, B1 => 
                           RF_RD2_DATA(19), B2 => n1816, ZN => n983);
   U2884 : XNOR2_X1 port map( A => n1889, B => 
                           DATAPATH_IxThird_stxALU_IN1_19_port, ZN => n576);
   U2885 : AOI21_X1 port map( B1 => n1957, B2 => n1886, A => n1955, ZN => n548)
                           ;
   U2886 : AOI22_X1 port map( A1 => n1909, A2 => n1798, B1 => 
                           DATAPATH_IxThird_stxALU1xN212, B2 => n1959, ZN => 
                           n550);
   U2887 : NOR2_X1 port map( A1 => n546, A2 => n1886, ZN => n544);
   U2888 : NAND2_X1 port map( A1 => n546, A2 => n1671, ZN => n540);
   U2889 : XNOR2_X1 port map( A => n1926, B => n1798, ZN => n553);
   U2890 : XNOR2_X1 port map( A => n2142, B => 
                           DATAPATH_IxThird_stxALU_IN1_21_port, ZN => n551);
   U2891 : OAI221_X1 port map( B1 => n1861, B2 => n1618, C1 => n1440, C2 => 
                           n1950, A => n997, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_21_port);
   U2892 : AOI22_X1 port map( A1 => RF_WR_DATAx17x, A2 => n1949, B1 => 
                           RF_RD1_DATA(17), B2 => n1888, ZN => n1007);
   U2893 : AOI22_X1 port map( A1 => RF_WR_DATAx20x, A2 => n1948, B1 => 
                           RF_RD1_DATA(20), B2 => n979, ZN => n994);
   U2894 : AOI22_X1 port map( A1 => RF_WR_DATAx18x, A2 => n1949, B1 => 
                           RF_RD1_DATA(18), B2 => n979, ZN => n1004);
   U2895 : AOI22_X1 port map( A1 => RF_WR_DATAx22x, A2 => n1949, B1 => 
                           RF_RD1_DATA(22), B2 => n1890, ZN => n988);
   U2896 : AOI22_X1 port map( A1 => RF_WR_DATAx30x, A2 => n1949, B1 => 
                           RF_RD1_DATA(30), B2 => n979, ZN => n1010);
   U2897 : AOI22_X1 port map( A1 => RF_WR_DATAx23x, A2 => n1949, B1 => 
                           RF_RD1_DATA(23), B2 => n1884, ZN => n1000);
   U2898 : AOI22_X1 port map( A1 => RF_WR_DATAx21x, A2 => n1948, B1 => 
                           RF_RD1_DATA(21), B2 => n979, ZN => n997);
   U2899 : XNOR2_X1 port map( A => n2147, B => 
                           DATAPATH_IxThird_stxALU_IN1_16_port, ZN => n618);
   U2900 : INV_X1 port map( A => n788, ZN => n2147);
   U2901 : AOI22_X1 port map( A1 => RF_WR_DATAx16x, A2 => n1949, B1 => 
                           RF_RD1_DATA(16), B2 => n1891, ZN => n991);
   U2902 : AOI21_X1 port map( B1 => n932, B2 => n931, A => n933, ZN => n929);
   U2903 : OAI21_X1 port map( B1 => n934, B2 => n791, A => n2196, ZN => n932);
   U2904 : AOI21_X1 port map( B1 => n282, B2 => n284, A => n815, ZN => n959);
   U2905 : OAI221_X1 port map( B1 => n1861, B2 => n1619, C1 => n1422, C2 => 
                           n1823, A => n1083, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_3_port);
   U2906 : OAI221_X1 port map( B1 => n1860, B2 => n1620, C1 => n1425, C2 => 
                           n1823, A => n1077, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_6_port);
   U2907 : OAI221_X1 port map( B1 => n1871, B2 => n1621, C1 => n1421, C2 => 
                           n1823, A => n1080, ZN => 
                           DATAPATH_IxThird_stxALU_IN1_2_port);
   U2908 : AOI21_X1 port map( B1 => n1775, B2 => n280, A => n2089, ZN => n1296)
                           ;
   U2909 : AOI22_X1 port map( A1 => n643, A2 => n1778, B1 => n2117, B2 => n644,
                           ZN => n638);
   U2910 : AOI22_X1 port map( A1 => n625, A2 => n1778, B1 => n2117, B2 => n628,
                           ZN => n620);
   U2911 : AOI22_X1 port map( A1 => n428, A2 => n1851, B1 => n2101, B2 => n431,
                           ZN => n423);
   U2912 : AOI22_X1 port map( A1 => n489, A2 => n1846, B1 => n2105, B2 => n490,
                           ZN => n483);
   U2913 : AOI22_X1 port map( A1 => n470, A2 => n1846, B1 => n2105, B2 => n473,
                           ZN => n465);
   U2914 : XNOR2_X1 port map( A => n394, B => n1840, ZN => n391);
   U2915 : XNOR2_X1 port map( A => n1846, B => n513, ZN => n510);
   U2916 : XNOR2_X1 port map( A => n1867, B => n348, ZN => n345);
   U2917 : XNOR2_X1 port map( A => n1852, B => n561, ZN => n558);
   U2918 : AOI22_X1 port map( A1 => n537, A2 => n1852, B1 => n2109, B2 => n538,
                           ZN => n532);
   U2919 : AOI22_X1 port map( A1 => n519, A2 => n1852, B1 => n2109, B2 => n522,
                           ZN => n514);
   U2920 : AOI22_X1 port map( A1 => n2125, A2 => n373, B1 => n374, B2 => n1840,
                           ZN => n367);
   U2921 : AOI22_X1 port map( A1 => n2125, A2 => n355, B1 => n356, B2 => n1840,
                           ZN => n349);
   U2922 : AOI22_X1 port map( A1 => n2121, A2 => n687, B1 => n688, B2 => n1867,
                           ZN => n682);
   U2923 : AOI22_X1 port map( A1 => n2121, A2 => n671, B1 => n672, B2 => n1867,
                           ZN => n665);
   U2924 : AOI21_X1 port map( B1 => n710, B2 => n1851, A => n1605, ZN => n702);
   U2925 : INV_X1 port map( A => n1867, ZN => n2121);
   U2926 : AOI222_X1 port map( A1 => DATAPATH_IxThird_stxALU1xN191, A2 => n1960
                           , B1 => n571, B2 => n1768, C1 => n1910, C2 => n1709,
                           ZN => n699);
   U2927 : OAI21_X1 port map( B1 => n455, B2 => n1851, A => n2098, ZN => n453);
   U2928 : OAI21_X1 port map( B1 => n337, B2 => n1867, A => n2120, ZN => n335);
   U2929 : INV_X1 port map( A => n1840, ZN => n2125);
   U2930 : INV_X1 port map( A => n1846, ZN => n2105);
   U2931 : INV_X1 port map( A => n1852, ZN => n2109);
   U2932 : AOI21_X1 port map( B1 => n543, B2 => n1852, A => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n555);
   U2933 : AOI21_X1 port map( B1 => n495, B2 => n1846, A => n1785, ZN => n507);
   U2934 : AOI21_X1 port map( B1 => n1867, B2 => n337, A => n1809, ZN => n340);
   U2935 : OAI22_X1 port map( A1 => n2101, A2 => n725, B1 => n726, B2 => n1851,
                           ZN => n420);
   U2936 : INV_X1 port map( A => n1839, ZN => n2101);
   U2937 : AOI22_X1 port map( A1 => n429, A2 => n2100, B1 => n457, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, ZN => n722);
   U2938 : AOI22_X1 port map( A1 => n471, A2 => n513, B1 => n495, B2 => n1785, 
                           ZN => n740);
   U2939 : AOI22_X1 port map( A1 => n520, A2 => n561, B1 => n543, B2 => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, ZN => n748);
   U2940 : INV_X1 port map( A => n1778, ZN => n2117);
   U2941 : AOI22_X1 port map( A1 => n338, A2 => n348, B1 => n337, B2 => n1809, 
                           ZN => n769);
   U2942 : AOI21_X1 port map( B1 => n357, B2 => n394, A => n2124, ZN => n776);
   U2943 : AOI21_X1 port map( B1 => n871, B2 => n870, A => n872, ZN => n868);
   U2944 : NAND2_X1 port map( A1 => n1241, A2 => n283, ZN => n284);
   U2945 : AOI21_X1 port map( B1 => n1591, B2 => n1735, A => n1748, ZN => n817)
                           ;
   U2946 : XNOR2_X1 port map( A => n1812, B => n1159, ZN => n1104);
   U2947 : AOI21_X1 port map( B1 => n906, B2 => n905, A => n907, ZN => n903);
   U2948 : INV_X1 port map( A => DATAPATH_IxThird_stxALU1xN222, ZN => n1979);
   U2949 : OAI22_X1 port map( A1 => n1979, A2 => n715, B1 => n716, B2 => n717, 
                           ZN => n708);
   U2950 : OAI21_X1 port map( B1 => n2077, B2 => n909, A => n910, ZN => n906);
   U2951 : XNOR2_X1 port map( A => n1878, B => n1145, ZN => n1103);
   U2952 : NAND2_X1 port map( A1 => CU_Ixcw2_i_10_port, A2 => n1750, ZN => 
                           n1451);
   U2953 : OAI221_X1 port map( B1 => n1861, B2 => n1622, C1 => n1450, C2 => 
                           n1950, A => n1013, ZN => 
                           DATAPATH_IxThird_stxALU1xN222);
   U2954 : OAI211_X1 port map( C1 => n1357, C2 => n1386, A => n850, B => n851, 
                           ZN => n835);
   U2955 : AOI22_X1 port map( A1 => RF_WR_DATAx1x, A2 => n1949, B1 => 
                           RF_RD1_DATA(1), B2 => n1947, ZN => n1086);
   U2956 : AOI22_X1 port map( A1 => RF_WR_DATAx9x, A2 => n1949, B1 => 
                           RF_RD1_DATA(9), B2 => n1946, ZN => n1040);
   U2957 : AOI22_X1 port map( A1 => RF_WR_DATAx8x, A2 => n1949, B1 => 
                           RF_RD1_DATA(8), B2 => n1947, ZN => n1037);
   U2958 : AOI22_X1 port map( A1 => RF_WR_DATAx28x, A2 => n1949, B1 => 
                           RF_RD1_DATA(28), B2 => n1890, ZN => n1029);
   U2959 : AOI22_X1 port map( A1 => RF_WR_DATAx15x, A2 => n1948, B1 => 
                           RF_RD1_DATA(15), B2 => n1884, ZN => n1046);
   U2960 : AOI22_X1 port map( A1 => RF_WR_DATAx11x, A2 => n1948, B1 => 
                           RF_RD1_DATA(11), B2 => n1888, ZN => n1057);
   U2961 : AOI22_X1 port map( A1 => RF_WR_DATAx14x, A2 => n1949, B1 => 
                           RF_RD1_DATA(14), B2 => n979, ZN => n1043);
   U2962 : AOI22_X1 port map( A1 => RF_WR_DATAx27x, A2 => n1949, B1 => 
                           RF_RD1_DATA(27), B2 => n1891, ZN => n1026);
   U2963 : AOI22_X1 port map( A1 => RF_WR_DATAx25x, A2 => n1949, B1 => 
                           RF_RD1_DATA(25), B2 => n1890, ZN => n1016);
   U2964 : AOI22_X1 port map( A1 => RF_WR_DATAx24x, A2 => n1949, B1 => 
                           RF_RD1_DATA(24), B2 => n1888, ZN => n1019);
   U2965 : AOI22_X1 port map( A1 => RF_WR_DATAx26x, A2 => n1949, B1 => 
                           RF_RD1_DATA(26), B2 => n1884, ZN => n1023);
   U2966 : AOI22_X1 port map( A1 => RF_WR_DATAx31x, A2 => n1949, B1 => 
                           RF_RD1_DATA(31), B2 => n1884, ZN => n1013);
   U2967 : NAND2_X1 port map( A1 => n1088, A2 => n1090, ZN => n976);
   U2968 : OAI21_X1 port map( B1 => n1820, B2 => n1592, A => n1775, ZN => n49);
   U2969 : OAI22_X1 port map( A1 => n1711, A2 => n818, B1 => n1760, B2 => n820,
                           ZN => DATAPATH_IxSecond_stxjump_target_31_port);
   U2970 : OAI22_X1 port map( A1 => n1711, A2 => n827, B1 => n828, B2 => n1760,
                           ZN => DATAPATH_IxSecond_stxjump_target_30_port);
   U2971 : INV_X1 port map( A => n817, ZN => n2087);
   U2972 : OAI21_X1 port map( B1 => n1824, B2 => n2158, A => n2041, ZN => n296)
                           ;
   U2973 : OAI21_X1 port map( B1 => n2158, B2 => n1824, A => n1212, ZN => n292)
                           ;
   U2974 : NAND2_X1 port map( A1 => n1829, A2 => n284, ZN => n282);
   U2975 : NAND2_X1 port map( A1 => n286, A2 => n1592, ZN => n279);
   U2976 : NAND4_X1 port map( A1 => n1654, A2 => n1581, A3 => n968, A4 => n967,
                           ZN => n294);
   U2977 : NOR2_X1 port map( A1 => n1198, A2 => n291, ZN => CU_Ixcw2_0_port);
   U2978 : NOR2_X1 port map( A1 => n1199, A2 => n291, ZN => CU_Ixcw2_1_port);
   U2979 : NOR2_X1 port map( A1 => n1200, A2 => n291, ZN => CU_Ixcw2_2_port);
   U2980 : NOR2_X1 port map( A1 => n1201, A2 => n291, ZN => CU_Ixcw2_3_port);
   U2981 : NOR2_X1 port map( A1 => n1202, A2 => n291, ZN => CU_Ixcw2_4_port);
   U2982 : NOR2_X1 port map( A1 => n1203, A2 => n291, ZN => CU_Ixcw2_5_port);
   U2983 : NOR2_X1 port map( A1 => n1204, A2 => n291, ZN => CU_Ixcw2_6_port);
   U2984 : OAI22_X1 port map( A1 => n795, A2 => n1729, B1 => n268, B2 => n797, 
                           ZN => DATAPATH_IxSecond_stxjump_target_7_port);
   U2985 : OAI22_X1 port map( A1 => n2053, A2 => n857, B1 => n1858, B2 => n858,
                           ZN => DATAPATH_IxSecond_stxjump_target_23_port);
   U2986 : OAI22_X1 port map( A1 => n2083, A2 => n938, B1 => n939, B2 => n1848,
                           ZN => DATAPATH_IxSecond_stxjump_target_11_port);
   U2987 : OAI22_X1 port map( A1 => n2057, A2 => n840, B1 => n1708, B2 => n841,
                           ZN => DATAPATH_IxSecond_stxjump_target_27_port);
   U2988 : OAI22_X1 port map( A1 => n2057, A2 => n846, B1 => n847, B2 => n1708,
                           ZN => DATAPATH_IxSecond_stxjump_target_26_port);
   U2989 : OAI21_X1 port map( B1 => n878, B2 => n2075, A => n1857, ZN => n901);
   U2990 : OAI22_X1 port map( A1 => n1729, A2 => n806, B1 => n268, B2 => n807, 
                           ZN => DATAPATH_IxSecond_stxjump_target_6_port);
   U2991 : OAI22_X1 port map( A1 => n1892, A2 => n918, B1 => n1841, B2 => n920,
                           ZN => DATAPATH_IxSecond_stxjump_target_14_port);
   U2992 : OAI22_X1 port map( A1 => n2065, A2 => n889, B1 => n1857, B2 => n890,
                           ZN => DATAPATH_IxSecond_stxjump_target_18_port);
   U2993 : OAI22_X1 port map( A1 => n2083, A2 => n947, B1 => n948, B2 => n1848,
                           ZN => DATAPATH_IxSecond_stxjump_target_10_port);
   U2994 : OAI22_X1 port map( A1 => n2053, A2 => n863, B1 => n864, B2 => n1858,
                           ZN => DATAPATH_IxSecond_stxjump_target_22_port);
   U2995 : OAI21_X1 port map( B1 => n1841, B2 => n921, A => n912, ZN => n925);
   U2996 : XNOR2_X1 port map( A => n927, B => n1841, ZN => 
                           DATAPATH_IxSecond_stxjump_target_12_port);
   U2997 : OAI21_X1 port map( B1 => n1917, B2 => n1859, A => n866, ZN => n865);
   U2998 : OAI211_X1 port map( C1 => n885, C2 => n1857, A => n886, B => n887, 
                           ZN => n884);
   U2999 : INV_X1 port map( A => n1848, ZN => n2083);
   U3000 : INV_X1 port map( A => n1857, ZN => n2065);
   U3001 : INV_X1 port map( A => n1858, ZN => n2053);
   U3002 : OR3_X1 port map( A1 => n291, A2 => n1205, A3 => n2093, ZN => n962);
   U3003 : INV_X1 port map( A => n1875, ZN => n2057);
   U3004 : OAI21_X1 port map( B1 => n1205, B2 => n291, A => n1451, ZN => n961);
   U3005 : NOR2_X1 port map( A1 => n1206, A2 => n291, ZN => RF_RD1_EN);
   U3006 : NOR2_X1 port map( A1 => n1207, A2 => n291, ZN => RF_RD2_EN);
   U3007 : NOR3_X1 port map( A1 => n2096, A2 => n1211, A3 => n291, ZN => n159);
   U3008 : AOI21_X1 port map( B1 => n876, B2 => n877, A => n878, ZN => n873);
   U3009 : OAI211_X1 port map( C1 => n1374, C2 => n1726, A => n2076, B => n1352
                           , ZN => n887);
   U3010 : OAI21_X1 port map( B1 => n291, B2 => n1211, A => n292, ZN => n165);
   U3011 : OAI211_X1 port map( C1 => n1373, C2 => n1726, A => n2076, B => n1351
                           , ZN => n894);
   U3012 : OAI211_X1 port map( C1 => n1372, C2 => n1726, A => n2076, B => n1350
                           , ZN => n877);
   U3013 : INV_X1 port map( A => n919, ZN => n2077);
   U3014 : OAI211_X1 port map( C1 => n1726, C2 => n1634, A => n2076, B => n1347
                           , ZN => n912);
   U3015 : OAI211_X1 port map( C1 => n1726, C2 => n1635, A => n2076, B => n1348
                           , ZN => n911);
   U3016 : AOI21_X1 port map( B1 => n936, B2 => n244, A => n794, ZN => n934);
   U3017 : AOI22_X1 port map( A1 => n1726, A2 => n1366, B1 => n1764, B2 => 
                           n1376, ZN => n945);
   U3018 : OAI22_X1 port map( A1 => n1370, A2 => n1764, B1 => n1380, B2 => 
                           n1771, ZN => n956);
   U3019 : AOI22_X1 port map( A1 => n1771, A2 => n1369, B1 => n1763, B2 => 
                           n1379, ZN => n958);
   U3020 : AOI22_X1 port map( A1 => n897, A2 => n1367, B1 => n1772, B2 => n1377
                           , ZN => n286);
   U3021 : INV_X1 port map( A => n1985, ZN => n1983);
   U3022 : INV_X1 port map( A => n1985, ZN => n1984);
   U3023 : INV_X1 port map( A => n1995, ZN => n1992);
   U3024 : INV_X1 port map( A => Rst, ZN => n1993);
   U3025 : INV_X1 port map( A => Rst, ZN => n1994);
   U3026 : INV_X1 port map( A => Rst, ZN => n1995);
   U3027 : NOR2_X1 port map( A1 => n1999, A2 => n2000, ZN => n1998);
   U3028 : OAI22_X1 port map( A1 => CU_IxN25, A2 => n2001, B1 => CU_IxN24, B2 
                           => n1998, ZN => CU_Ixcw_LUT_0_port);
   U3029 : AOI21_X1 port map( B1 => CU_IxN23, B2 => n1999, A => n2001, ZN => 
                           n1996);
   U3030 : NOR2_X1 port map( A1 => n1998, A2 => n1996, ZN => CU_Ixcw_LUT_1_port
                           );
   U3031 : NOR3_X1 port map( A1 => n2001, A2 => CU_IxN25, A3 => CU_IxN23, ZN =>
                           CU_Ixcw_LUT_2_port);
   U3032 : NOR3_X1 port map( A1 => n2001, A2 => CU_IxN23, A3 => n1999, ZN => 
                           CU_Ixcw_LUT_4_port);
   U3033 : OAI21_X1 port map( B1 => CU_IxN24, B2 => n2000, A => CU_IxN25, ZN =>
                           CU_Ixcw_LUT_5_port);
   U3034 : AOI21_X1 port map( B1 => CU_IxN24, B2 => CU_IxN23, A => n1999, ZN =>
                           CU_Ixcw_LUT_7_port);
   U3035 : OAI22_X1 port map( A1 => CU_IxN24, A2 => n1999, B1 => n1998, B2 => 
                           n2001, ZN => CU_Ixcw_LUT_8_port);
   U3036 : NOR2_X1 port map( A1 => CU_IxN24, A2 => CU_IxN25, ZN => 
                           CU_Ixcw_LUT_10_port);
   U3037 : NAND2_X1 port map( A1 => CU_Ixcw_LUT_10_port, A2 => CU_IxN23, ZN => 
                           n1997);
   U3038 : OAI21_X1 port map( B1 => n1999, B2 => n2001, A => n1997, ZN => 
                           CU_Ixcw_LUT_15_port);
   U3039 : NAND2_X1 port map( A1 => CU_IxN24, A2 => n1998, ZN => 
                           CU_Ixcw_LUT_16_port);
   U3040 : AND2_X1 port map( A1 => n2001, A2 => n1998, ZN => CU_Ixcw_LUT_9_port
                           );
   U3041 : MUX2_X1 port map( A => n1716, B => 
                           DATAPATH_IxThird_stxALU_IN1_1_port, S => n1990, Z =>
                           n2210);
   U3042 : MUX2_X1 port map( A => n1734, B => 
                           DATAPATH_IxThird_stxALU_IN1_3_port, S => n1990, Z =>
                           n2306);
   U3043 : MUX2_X1 port map( A => n2210, B => n2306, S => n1989, Z => n2211);
   U3044 : MUX2_X1 port map( A => n1791, B => 
                           DATAPATH_IxThird_stxALU_IN1_5_port, S => n1990, Z =>
                           n2305);
   U3045 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_6_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_7_port, S => n1990, Z =>
                           n2308);
   U3046 : MUX2_X1 port map( A => n2305, B => n2308, S => n1989, Z => n2328);
   U3047 : MUX2_X1 port map( A => n2211, B => n2328, S => n1681, Z => n2212);
   U3048 : MUX2_X1 port map( A => n1809, B => n1794, S => n1990, Z => n2307);
   U3049 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_10_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_11_port, S => n1990, Z 
                           => n2216);
   U3050 : MUX2_X1 port map( A => n2307, B => n2216, S => n1989, Z => n2327);
   U3051 : MUX2_X1 port map( A => n1796, B => 
                           DATAPATH_IxThird_stxALU_IN1_13_port, S => n1990, Z 
                           => n2215);
   U3052 : MUX2_X1 port map( A => n1787, B => n1797, S => n1990, Z => n2218);
   U3053 : MUX2_X1 port map( A => n2215, B => n2218, S => n1989, Z => n2231);
   U3054 : MUX2_X1 port map( A => n2327, B => n2231, S => n1681, Z => n2356);
   U3055 : MUX2_X1 port map( A => n2212, B => n2356, S => n1987, Z => n2213);
   U3056 : MUX2_X1 port map( A => n1655, B => n1668, S => n1990, Z => n2217);
   U3057 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_18_port, B => 
                           n1663, S => n1990, Z => n2220);
   U3058 : MUX2_X1 port map( A => n2217, B => n2220, S => n1989, Z => n2230);
   U3059 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_20_port, B => 
                           n1886, S => n1990, Z => n2219);
   U3060 : MUX2_X1 port map( A => n1670, B => n1784, S => n1990, Z => n2222);
   U3061 : MUX2_X1 port map( A => n2219, B => n2222, S => n1989, Z => n2233);
   U3062 : MUX2_X1 port map( A => n2230, B => n2233, S => n1681, Z => n2355);
   U3063 : MUX2_X1 port map( A => n1785, B => n1674, S => n1990, Z => n2221);
   U3064 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_26_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_27_port, S => n1990, Z 
                           => n2224);
   U3065 : MUX2_X1 port map( A => n2221, B => n2224, S => n1989, Z => n2232);
   U3066 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_28_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_29_port, S => n1990, Z 
                           => n2223);
   U3067 : MUX2_X1 port map( A => n1783, B => n1872, S => n1990, Z => n2225);
   U3068 : MUX2_X1 port map( A => n2223, B => n2225, S => n1989, Z => n2234);
   U3069 : MUX2_X1 port map( A => n2232, B => n2234, S => n1681, Z => n2293);
   U3070 : MUX2_X1 port map( A => n2355, B => n2293, S => n1987, Z => n2261);
   U3071 : MUX2_X1 port map( A => n2213, B => n2261, S => n1983, Z => n2214);
   U3072 : MUX2_X1 port map( A => n2214, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN191);
   U3073 : MUX2_X1 port map( A => n2216, B => n2215, S => n1989, Z => n2341);
   U3074 : MUX2_X1 port map( A => n2218, B => n2217, S => n1989, Z => n2249);
   U3075 : MUX2_X1 port map( A => n2341, B => n2249, S => n1681, Z => n2310);
   U3076 : MUX2_X1 port map( A => n2220, B => n2219, S => n1989, Z => n2248);
   U3077 : MUX2_X1 port map( A => n2222, B => n2221, S => n1989, Z => n2251);
   U3078 : MUX2_X1 port map( A => n2248, B => n2251, S => n1681, Z => n2269);
   U3079 : MUX2_X1 port map( A => n2310, B => n2269, S => n1987, Z => n2226);
   U3080 : MUX2_X1 port map( A => n2224, B => n2223, S => n1989, Z => n2250);
   U3081 : MUX2_X1 port map( A => n2225, B => n1873, S => n1989, Z => n2252);
   U3082 : MUX2_X1 port map( A => n2250, B => n2252, S => n1681, Z => n2268);
   U3083 : MUX2_X1 port map( A => n2268, B => n1873, S => n1987, Z => n2297);
   U3084 : MUX2_X1 port map( A => n2226, B => n2297, S => n1983, Z => n2227);
   U3085 : MUX2_X1 port map( A => n2227, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN201);
   U3086 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_11_port, B => 
                           n1796, S => n1990, Z => n2276);
   U3087 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_13_port, B => 
                           n1787, S => n1990, Z => n2238);
   U3088 : MUX2_X1 port map( A => n2276, B => n2238, S => n1989, Z => n2348);
   U3089 : MUX2_X1 port map( A => n1797, B => n1655, S => n1990, Z => n2237);
   U3090 : MUX2_X1 port map( A => n1669, B => 
                           DATAPATH_IxThird_stxALU_IN1_18_port, S => n1990, Z 
                           => n2240);
   U3091 : MUX2_X1 port map( A => n2237, B => n2240, S => n1989, Z => n2256);
   U3092 : MUX2_X1 port map( A => n2348, B => n2256, S => n1681, Z => n2322);
   U3093 : MUX2_X1 port map( A => n1663, B => 
                           DATAPATH_IxThird_stxALU_IN1_20_port, S => n1990, Z 
                           => n2239);
   U3094 : MUX2_X1 port map( A => n1671, B => n1670, S => n1990, Z => n2242);
   U3095 : MUX2_X1 port map( A => n2239, B => n2242, S => n1989, Z => n2255);
   U3096 : MUX2_X1 port map( A => n1784, B => n1785, S => n1990, Z => n2241);
   U3097 : MUX2_X1 port map( A => n1674, B => 
                           DATAPATH_IxThird_stxALU_IN1_26_port, S => n1990, Z 
                           => n2244);
   U3098 : MUX2_X1 port map( A => n2241, B => n2244, S => n1989, Z => n2258);
   U3099 : MUX2_X1 port map( A => n2255, B => n2258, S => n1681, Z => n2272);
   U3100 : MUX2_X1 port map( A => n2322, B => n2272, S => n1987, Z => n2228);
   U3101 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_27_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_28_port, S => n1990, Z 
                           => n2243);
   U3102 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_29_port, B => 
                           n1783, S => n1990, Z => n2245);
   U3103 : MUX2_X1 port map( A => n2243, B => n2245, S => n1989, Z => n2257);
   U3104 : MUX2_X1 port map( A => n2257, B => n1873, S => n1681, Z => n2271);
   U3105 : MUX2_X1 port map( A => n2271, B => n1873, S => n1987, Z => n2299);
   U3106 : MUX2_X1 port map( A => n2228, B => n2299, S => n1983, Z => n2229);
   U3107 : MUX2_X1 port map( A => n2229, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN202);
   U3108 : MUX2_X1 port map( A => n2231, B => n2230, S => n1681, Z => n2329);
   U3109 : MUX2_X1 port map( A => n2233, B => n2232, S => n1681, Z => n2283);
   U3110 : MUX2_X1 port map( A => n2329, B => n2283, S => n1987, Z => n2235);
   U3111 : MUX2_X1 port map( A => n2234, B => n1873, S => n1681, Z => n2282);
   U3112 : MUX2_X1 port map( A => n2282, B => n1873, S => n1987, Z => n2301);
   U3113 : MUX2_X1 port map( A => n2235, B => n2301, S => n1983, Z => n2236);
   U3114 : MUX2_X1 port map( A => n2236, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN203);
   U3115 : MUX2_X1 port map( A => n2238, B => n2237, S => n1989, Z => n2277);
   U3116 : MUX2_X1 port map( A => n2240, B => n2239, S => n1989, Z => n2264);
   U3117 : MUX2_X1 port map( A => n2277, B => n2264, S => n1681, Z => n2336);
   U3118 : MUX2_X1 port map( A => n2242, B => n2241, S => n1989, Z => n2263);
   U3119 : MUX2_X1 port map( A => n2244, B => n2243, S => n1989, Z => n2266);
   U3120 : MUX2_X1 port map( A => n2263, B => n2266, S => n1681, Z => n2286);
   U3121 : MUX2_X1 port map( A => n2336, B => n2286, S => n1987, Z => n2246);
   U3122 : MUX2_X1 port map( A => n2245, B => n1873, S => n1989, Z => n2265);
   U3123 : MUX2_X1 port map( A => n2265, B => n1873, S => n1681, Z => n2285);
   U3124 : MUX2_X1 port map( A => n2285, B => n1873, S => n1987, Z => n2303);
   U3125 : MUX2_X1 port map( A => n2246, B => n2303, S => n1983, Z => n2247);
   U3126 : MUX2_X1 port map( A => n2247, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN204);
   U3127 : MUX2_X1 port map( A => n2249, B => n2248, S => n1681, Z => n2343);
   U3128 : MUX2_X1 port map( A => n2251, B => n2250, S => n1681, Z => n2289);
   U3129 : MUX2_X1 port map( A => n2343, B => n2289, S => n1987, Z => n2253);
   U3130 : MUX2_X1 port map( A => n2252, B => n1873, S => n1681, Z => n2288);
   U3131 : MUX2_X1 port map( A => n2288, B => n1873, S => n1987, Z => n2315);
   U3132 : MUX2_X1 port map( A => n2253, B => n2315, S => n1983, Z => n2254);
   U3133 : MUX2_X1 port map( A => n2254, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN205);
   U3134 : MUX2_X1 port map( A => n2256, B => n2255, S => n1681, Z => n2350);
   U3135 : MUX2_X1 port map( A => n2258, B => n2257, S => n1681, Z => n2291);
   U3136 : MUX2_X1 port map( A => n2350, B => n2291, S => n1987, Z => n2259);
   U3137 : MUX2_X1 port map( A => n2259, B => n1873, S => n1983, Z => n2260);
   U3138 : MUX2_X1 port map( A => n2260, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN206);
   U3139 : MUX2_X1 port map( A => n2261, B => n1873, S => n1983, Z => n2262);
   U3140 : MUX2_X1 port map( A => n2262, B => n1873, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN207);
   U3141 : MUX2_X1 port map( A => n2264, B => n2263, S => n1681, Z => n2360);
   U3142 : MUX2_X1 port map( A => n2266, B => n2265, S => n1681, Z => n2295);
   U3143 : MUX2_X1 port map( A => n2360, B => n2295, S => n1987, Z => n2279);
   U3144 : MUX2_X1 port map( A => n2279, B => n1873, S => n1983, Z => n2267);
   U3145 : MUX2_X1 port map( A => n2267, B => n1874, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN208);
   U3146 : MUX2_X1 port map( A => n2269, B => n2268, S => n1987, Z => n2312);
   U3147 : MUX2_X1 port map( A => n2312, B => n1874, S => n1983, Z => n2270);
   U3148 : MUX2_X1 port map( A => n2270, B => n1874, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN209);
   U3149 : MUX2_X1 port map( A => n2272, B => n2271, S => n1987, Z => n2324);
   U3150 : MUX2_X1 port map( A => n2324, B => n1874, S => n1983, Z => n2273);
   U3151 : MUX2_X1 port map( A => n2273, B => n1874, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN210);
   U3152 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_1_port, B => 
                           n1734, S => n1990, Z => n2274);
   U3153 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_3_port, B => 
                           n1791, S => n1990, Z => n2318);
   U3154 : MUX2_X1 port map( A => n2274, B => n2318, S => n1989, Z => n2275);
   U3155 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_5_port, B => 
                           DATAPATH_IxThird_stxALU_IN1_6_port, S => n1990, Z =>
                           n2317);
   U3156 : MUX2_X1 port map( A => DATAPATH_IxThird_stxALU_IN1_7_port, B => 
                           n1809, S => n1990, Z => n2320);
   U3157 : MUX2_X1 port map( A => n2317, B => n2320, S => n1989, Z => n2335);
   U3158 : MUX2_X1 port map( A => n2275, B => n2335, S => n1681, Z => n2278);
   U3159 : MUX2_X1 port map( A => n1794, B => 
                           DATAPATH_IxThird_stxALU_IN1_10_port, S => n1990, Z 
                           => n2319);
   U3160 : MUX2_X1 port map( A => n2319, B => n2276, S => n1989, Z => n2334);
   U3161 : MUX2_X1 port map( A => n2334, B => n2277, S => n1681, Z => n2361);
   U3162 : MUX2_X1 port map( A => n2278, B => n2361, S => n1987, Z => n2280);
   U3163 : MUX2_X1 port map( A => n2280, B => n2279, S => n1983, Z => n2281);
   U3164 : MUX2_X1 port map( A => n2281, B => n1874, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN192);
   U3165 : MUX2_X1 port map( A => n2283, B => n2282, S => n1987, Z => n2331);
   U3166 : MUX2_X1 port map( A => n2331, B => n1874, S => n1984, Z => n2284);
   U3167 : MUX2_X1 port map( A => n2284, B => n1874, S => n1980, Z => 
                           DATAPATH_IxThird_stxALU1xN211);
   U3168 : MUX2_X1 port map( A => n2286, B => n2285, S => n1987, Z => n2338);
   U3169 : MUX2_X1 port map( A => n2338, B => n1874, S => n1984, Z => n2287);
   U3170 : MUX2_X1 port map( A => n2287, B => n1874, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN212);
   U3171 : MUX2_X1 port map( A => n2289, B => n2288, S => n1987, Z => n2345);
   U3172 : MUX2_X1 port map( A => n2345, B => n1873, S => n1984, Z => n2290);
   U3173 : MUX2_X1 port map( A => n2290, B => n1873, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN213);
   U3174 : MUX2_X1 port map( A => n2291, B => n1873, S => n1987, Z => n2352);
   U3175 : MUX2_X1 port map( A => n2352, B => n1873, S => n1984, Z => n2292);
   U3176 : MUX2_X1 port map( A => n2292, B => n1873, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN214);
   U3177 : MUX2_X1 port map( A => n2293, B => n1873, S => n1987, Z => n2357);
   U3178 : MUX2_X1 port map( A => n2357, B => n1872, S => n1984, Z => n2294);
   U3179 : MUX2_X1 port map( A => n2294, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN215);
   U3180 : MUX2_X1 port map( A => n2295, B => n1872, S => n1987, Z => n2362);
   U3181 : MUX2_X1 port map( A => n2362, B => n1872, S => n1984, Z => n2296);
   U3182 : MUX2_X1 port map( A => n2296, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN216);
   U3183 : MUX2_X1 port map( A => n2297, B => n1872, S => n1984, Z => n2298);
   U3184 : MUX2_X1 port map( A => n2298, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN217);
   U3185 : MUX2_X1 port map( A => n2299, B => n1872, S => n1984, Z => n2300);
   U3186 : MUX2_X1 port map( A => n2300, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN218);
   U3187 : MUX2_X1 port map( A => n2301, B => n1872, S => n1984, Z => n2302);
   U3188 : MUX2_X1 port map( A => n2302, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN219);
   U3189 : MUX2_X1 port map( A => n2303, B => n1872, S => n1984, Z => n2304);
   U3190 : MUX2_X1 port map( A => n2304, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN220);
   U3191 : MUX2_X1 port map( A => n2306, B => n2305, S => n1989, Z => n2309);
   U3192 : MUX2_X1 port map( A => n2308, B => n2307, S => n1989, Z => n2342);
   U3193 : MUX2_X1 port map( A => n2309, B => n2342, S => n1681, Z => n2311);
   U3194 : MUX2_X1 port map( A => n2311, B => n2310, S => n1987, Z => n2313);
   U3195 : MUX2_X1 port map( A => n2313, B => n2312, S => n1984, Z => n2314);
   U3196 : MUX2_X1 port map( A => n2314, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN193);
   U3197 : MUX2_X1 port map( A => n2315, B => n1872, S => n1984, Z => n2316);
   U3198 : MUX2_X1 port map( A => n2316, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN221);
   U3199 : MUX2_X1 port map( A => n2318, B => n2317, S => n1989, Z => n2321);
   U3200 : MUX2_X1 port map( A => n2320, B => n2319, S => n1989, Z => n2349);
   U3201 : MUX2_X1 port map( A => n2321, B => n2349, S => n1681, Z => n2323);
   U3202 : MUX2_X1 port map( A => n2323, B => n2322, S => n1987, Z => n2325);
   U3203 : MUX2_X1 port map( A => n2325, B => n2324, S => n1983, Z => n2326);
   U3204 : MUX2_X1 port map( A => n2326, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN194);
   U3205 : MUX2_X1 port map( A => n2328, B => n2327, S => n1681, Z => n2330);
   U3206 : MUX2_X1 port map( A => n2330, B => n2329, S => n1987, Z => n2332);
   U3207 : MUX2_X1 port map( A => n2332, B => n2331, S => n1983, Z => n2333);
   U3208 : MUX2_X1 port map( A => n2333, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN195);
   U3209 : MUX2_X1 port map( A => n2335, B => n2334, S => n1681, Z => n2337);
   U3210 : MUX2_X1 port map( A => n2337, B => n2336, S => n1987, Z => n2339);
   U3211 : MUX2_X1 port map( A => n2339, B => n2338, S => n1983, Z => n2340);
   U3212 : MUX2_X1 port map( A => n2340, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN196);
   U3213 : MUX2_X1 port map( A => n2342, B => n2341, S => n1681, Z => n2344);
   U3214 : MUX2_X1 port map( A => n2344, B => n2343, S => n1987, Z => n2346);
   U3215 : MUX2_X1 port map( A => n2346, B => n2345, S => n1984, Z => n2347);
   U3216 : MUX2_X1 port map( A => n2347, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN197);
   U3217 : MUX2_X1 port map( A => n2349, B => n2348, S => n1681, Z => n2351);
   U3218 : MUX2_X1 port map( A => n2351, B => n2350, S => n1987, Z => n2353);
   U3219 : MUX2_X1 port map( A => n2353, B => n2352, S => n1984, Z => n2354);
   U3220 : MUX2_X1 port map( A => n2354, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN198);
   U3221 : MUX2_X1 port map( A => n2356, B => n2355, S => n1987, Z => n2358);
   U3222 : MUX2_X1 port map( A => n2358, B => n2357, S => n1984, Z => n2359);
   U3223 : MUX2_X1 port map( A => n2359, B => n1872, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN199);
   U3224 : MUX2_X1 port map( A => n2361, B => n2360, S => n1987, Z => n2363);
   U3225 : MUX2_X1 port map( A => n2363, B => n2362, S => n1984, Z => n2364);
   U3226 : MUX2_X1 port map( A => n2364, B => n1874, S => n1981, Z => 
                           DATAPATH_IxThird_stxALU1xN200);

end SYN_RV32I_rtl;
