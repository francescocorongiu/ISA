
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RV32I is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RV32I;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RV32I.all;

entity RV32I is

   port( Clk, Rst : in std_logic;  IRAM_DOUT, RF_RD1_DATA, RF_RD2_DATA, 
         DRAM_DOUT : in std_logic_vector (31 downto 0);  IRAM_ADD : out 
         std_logic_vector (31 downto 0);  RF_RD1_EN, RF_RD2_EN, RF_WR_EN : out 
         std_logic;  RF_RD1_ADD, RF_RD2_ADD, RF_WR_ADD : out std_logic_vector 
         (4 downto 0);  RF_WR_DATA : out std_logic_vector (31 downto 0);  
         DRAM_WE, DRAM_RE : out std_logic;  DRAM_ADD, DRAM_DIN : out 
         std_logic_vector (31 downto 0));

end RV32I;

architecture SYN_RV32I_rtl of RV32I is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, CU_IxN53, CU_IxN52, 
      DATAPATH_IxWR_ADD_MEM_fu_0_port, DATAPATH_IxWR_ADD_MEM_fu_1_port, 
      DATAPATH_IxWR_ADD_MEM_fu_2_port, DATAPATH_IxWR_ADD_MEM_fu_3_port, 
      DATAPATH_IxWR_ADD_MEM_fu_4_port, DATAPATH_IxPC4_0_port, 
      DATAPATH_IxPC4_1_port, DATAPATH_IxINSTR_7_port, DATAPATH_IxINSTR_8_port, 
      DATAPATH_IxINSTR_9_port, DATAPATH_IxINSTR_10_port, 
      DATAPATH_IxINSTR_11_port, DATAPATH_IxSecond_stxWRADD_d1_0_port, 
      DATAPATH_IxSecond_stxWRADD_d1_1_port, 
      DATAPATH_IxSecond_stxWRADD_d1_2_port, 
      DATAPATH_IxSecond_stxWRADD_d1_3_port, 
      DATAPATH_IxSecond_stxWRADD_d1_4_port, 
      DATAPATH_IxThird_stxALU_out_i_0_port, 
      DATAPATH_IxThird_stxALU_out_i_1_port, 
      DATAPATH_IxThird_stxALU_out_i_2_port, 
      DATAPATH_IxThird_stxALU_out_i_3_port, 
      DATAPATH_IxThird_stxALU_out_i_4_port, 
      DATAPATH_IxThird_stxALU_out_i_5_port, 
      DATAPATH_IxThird_stxALU_out_i_6_port, 
      DATAPATH_IxThird_stxALU_out_i_7_port, 
      DATAPATH_IxThird_stxALU_out_i_8_port, 
      DATAPATH_IxThird_stxALU_out_i_9_port, 
      DATAPATH_IxThird_stxALU_out_i_10_port, 
      DATAPATH_IxThird_stxALU_out_i_11_port, 
      DATAPATH_IxThird_stxALU_out_i_12_port, 
      DATAPATH_IxThird_stxALU_out_i_13_port, 
      DATAPATH_IxThird_stxALU_out_i_14_port, 
      DATAPATH_IxThird_stxALU_out_i_15_port, 
      DATAPATH_IxThird_stxALU_out_i_16_port, 
      DATAPATH_IxThird_stxALU_out_i_17_port, 
      DATAPATH_IxThird_stxALU_out_i_18_port, 
      DATAPATH_IxThird_stxALU_out_i_19_port, 
      DATAPATH_IxThird_stxALU_out_i_20_port, 
      DATAPATH_IxThird_stxALU_out_i_21_port, 
      DATAPATH_IxThird_stxALU_out_i_22_port, 
      DATAPATH_IxThird_stxALU_out_i_23_port, 
      DATAPATH_IxThird_stxALU_out_i_24_port, 
      DATAPATH_IxThird_stxALU_out_i_25_port, 
      DATAPATH_IxThird_stxALU_out_i_26_port, 
      DATAPATH_IxThird_stxALU_out_i_27_port, 
      DATAPATH_IxThird_stxALU_out_i_28_port, 
      DATAPATH_IxThird_stxALU_out_i_29_port, 
      DATAPATH_IxThird_stxALU_out_i_30_port, 
      DATAPATH_IxThird_stxALU_out_i_31_port, DATAPATH_IxThird_stxALU1xN297, 
      DATAPATH_IxThird_stxALU1xN296, DATAPATH_IxThird_stxALU1xN295, 
      DATAPATH_IxThird_stxALU1xN294, DATAPATH_IxThird_stxALU1xN293, 
      DATAPATH_IxThird_stxALU1xN292, DATAPATH_IxThird_stxALU1xN291, 
      DATAPATH_IxThird_stxALU1xN290, DATAPATH_IxThird_stxALU1xN289, 
      DATAPATH_IxThird_stxALU1xN288, DATAPATH_IxThird_stxALU1xN287, 
      DATAPATH_IxThird_stxALU1xN286, DATAPATH_IxThird_stxALU1xN285, 
      DATAPATH_IxThird_stxALU1xN284, DATAPATH_IxThird_stxALU1xN283, 
      DATAPATH_IxThird_stxALU1xN282, DATAPATH_IxThird_stxALU1xN281, 
      DATAPATH_IxThird_stxALU1xN280, DATAPATH_IxThird_stxALU1xN279, 
      DATAPATH_IxThird_stxALU1xN278, DATAPATH_IxThird_stxALU1xN277, 
      DATAPATH_IxThird_stxALU1xN276, DATAPATH_IxThird_stxALU1xN275, 
      DATAPATH_IxThird_stxALU1xN274, DATAPATH_IxThird_stxALU1xN273, 
      DATAPATH_IxThird_stxALU1xN272, DATAPATH_IxThird_stxALU1xN271, 
      DATAPATH_IxThird_stxALU1xN270, DATAPATH_IxThird_stxALU1xN269, 
      DATAPATH_IxThird_stxALU1xN268, DATAPATH_IxThird_stxALU1xN267, n21, n23, 
      n24, n26, n27, n28, n29, n33, n35, n36, n37, n38, n41, n45, n47, n63, n64
      , n65, n68, n70, n72, n73, n74, n76, n78, n79, n81, n82, n83, n86, n87, 
      n89, n90, n91, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104, 
      n106, n109, n110, n111, n112, n114, n117, n118, n120, n121, n122, n125, 
      n126, n128, n129, n130, n133, n134, n136, n137, n138, n141, n142, n144, 
      n145, n146, n149, n150, n152, n153, n154, n157, n158, n160, n161, n162, 
      n165, n166, n168, n169, n170, n171, n172, n176, n177, n179, n181, n182, 
      n184, n185, n186, n187, n188, n189, n191, n196, n198, n199, n200, n203, 
      n204, n205, n206, n207, n208, n211, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230, n231, 
      n232, n233, n234, n235, n236, n237, n239, n240, n241, n242, n243, n244, 
      n245, n247, n249, n250, n251, n252, n254, n255, n256, n257, n259, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n274, 
      n275, n276, n278, n279, n280, n281, n283, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n295, n296, n297, n298, n299, n300, n301, n302, 
      n304, n305, n306, n307, n308, n309, n310, n311, n314, n315, n317, n318, 
      n319, n320, n321, n322, n323, n325, n326, n327, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n352, n353, n354, n355, n356, n357, n358, 
      n361, n362, n364, n365, n366, n367, n368, n369, n370, n372, n373, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n390, n391, n392, n393, n394, n395, n398, n399, n400, n402, n403, 
      n404, n405, n406, n407, n408, n411, n412, n414, n415, n416, n417, n418, 
      n419, n420, n422, n423, n424, n425, n426, n428, n429, n430, n431, n433, 
      n435, n436, n437, n439, n441, n442, n444, n445, n446, n447, n449, n450, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n462, n463, n464, 
      n465, n466, n467, n468, n471, n472, n474, n475, n476, n477, n478, n479, 
      n480, n482, n483, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n500, n501, n502, n503, n504, n505, n506, 
      n507, n509, n510, n511, n512, n513, n514, n515, n518, n519, n521, n522, 
      n523, n524, n525, n526, n527, n529, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n558, n560, n561, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n617, n618, n620, n621, n622, n623, n624, n626, n627, n628, n629, n630, 
      n631, n632, n634, n635, n637, n638, n639, n640, n641, n643, n644, n645, 
      n647, n648, n649, n651, n652, n654, n655, n656, n658, n659, n662, n663, 
      n665, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, 
      n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, 
      n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, 
      n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, 
      n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
      n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
      n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, 
      n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, 
      n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
      n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
      n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, 
      n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, 
      n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, 
      n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
      n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116 : std_logic;

begin
   IRAM_ADD <= ( IRAM_ADD_31_port, IRAM_ADD_30_port, IRAM_ADD_29_port, 
      IRAM_ADD_28_port, IRAM_ADD_27_port, IRAM_ADD_26_port, IRAM_ADD_25_port, 
      IRAM_ADD_24_port, IRAM_ADD_23_port, IRAM_ADD_22_port, IRAM_ADD_21_port, 
      IRAM_ADD_20_port, IRAM_ADD_19_port, IRAM_ADD_18_port, IRAM_ADD_17_port, 
      IRAM_ADD_16_port, IRAM_ADD_15_port, IRAM_ADD_14_port, IRAM_ADD_13_port, 
      IRAM_ADD_12_port, IRAM_ADD_11_port, IRAM_ADD_10_port, IRAM_ADD_9_port, 
      IRAM_ADD_8_port, IRAM_ADD_7_port, IRAM_ADD_6_port, IRAM_ADD_5_port, 
      IRAM_ADD_4_port, IRAM_ADD_3_port, IRAM_ADD_2_port, DATAPATH_IxPC4_1_port,
      DATAPATH_IxPC4_0_port );
   
   CU_Ixstate_var_regx0x : DFFR_X1 port map( D => CU_IxN52, CK => Clk, RN => 
                           Rst, Q => n_1000, QN => n698);
   DATAPATH_IxThird_stxB_FORWARD_out_regx0x : DFF_X1 port map( D => n823, CK =>
                           Clk, Q => DRAM_DIN(0), QN => n_1001);
   DATAPATH_IxThird_stxB_FORWARD_out_regx1x : DFF_X1 port map( D => n821, CK =>
                           Clk, Q => DRAM_DIN(1), QN => n_1002);
   DATAPATH_IxThird_stxB_FORWARD_out_regx2x : DFF_X1 port map( D => n819, CK =>
                           Clk, Q => DRAM_DIN(2), QN => n_1003);
   DATAPATH_IxThird_stxB_FORWARD_out_regx3x : DFF_X1 port map( D => n817, CK =>
                           Clk, Q => DRAM_DIN(3), QN => n_1004);
   DATAPATH_IxThird_stxB_FORWARD_out_regx4x : DFF_X1 port map( D => 
                           RF_RD2_DATA(4), CK => Clk, Q => DRAM_DIN(4), QN => 
                           n_1005);
   DATAPATH_IxThird_stxB_FORWARD_out_regx5x : DFF_X1 port map( D => 
                           RF_RD2_DATA(5), CK => Clk, Q => DRAM_DIN(5), QN => 
                           n_1006);
   DATAPATH_IxThird_stxB_FORWARD_out_regx6x : DFF_X1 port map( D => 
                           RF_RD2_DATA(6), CK => Clk, Q => DRAM_DIN(6), QN => 
                           n_1007);
   DATAPATH_IxThird_stxB_FORWARD_out_regx7x : DFF_X1 port map( D => 
                           RF_RD2_DATA(7), CK => Clk, Q => DRAM_DIN(7), QN => 
                           n_1008);
   DATAPATH_IxThird_stxB_FORWARD_out_regx8x : DFF_X1 port map( D => 
                           RF_RD2_DATA(8), CK => Clk, Q => DRAM_DIN(8), QN => 
                           n_1009);
   DATAPATH_IxThird_stxB_FORWARD_out_regx9x : DFF_X1 port map( D => 
                           RF_RD2_DATA(9), CK => Clk, Q => DRAM_DIN(9), QN => 
                           n_1010);
   DATAPATH_IxThird_stxB_FORWARD_out_regx10x : DFF_X1 port map( D => 
                           RF_RD2_DATA(10), CK => Clk, Q => DRAM_DIN(10), QN =>
                           n_1011);
   DATAPATH_IxThird_stxB_FORWARD_out_regx11x : DFF_X1 port map( D => 
                           RF_RD2_DATA(11), CK => Clk, Q => DRAM_DIN(11), QN =>
                           n_1012);
   DATAPATH_IxThird_stxB_FORWARD_out_regx12x : DFF_X1 port map( D => 
                           RF_RD2_DATA(12), CK => Clk, Q => DRAM_DIN(12), QN =>
                           n_1013);
   DATAPATH_IxThird_stxB_FORWARD_out_regx13x : DFF_X1 port map( D => 
                           RF_RD2_DATA(13), CK => Clk, Q => DRAM_DIN(13), QN =>
                           n_1014);
   DATAPATH_IxThird_stxB_FORWARD_out_regx14x : DFF_X1 port map( D => 
                           RF_RD2_DATA(14), CK => Clk, Q => DRAM_DIN(14), QN =>
                           n_1015);
   DATAPATH_IxThird_stxB_FORWARD_out_regx15x : DFF_X1 port map( D => 
                           RF_RD2_DATA(15), CK => Clk, Q => DRAM_DIN(15), QN =>
                           n_1016);
   DATAPATH_IxThird_stxB_FORWARD_out_regx16x : DFF_X1 port map( D => 
                           RF_RD2_DATA(16), CK => Clk, Q => DRAM_DIN(16), QN =>
                           n_1017);
   DATAPATH_IxThird_stxB_FORWARD_out_regx17x : DFF_X1 port map( D => 
                           RF_RD2_DATA(17), CK => Clk, Q => DRAM_DIN(17), QN =>
                           n_1018);
   DATAPATH_IxThird_stxB_FORWARD_out_regx18x : DFF_X1 port map( D => 
                           RF_RD2_DATA(18), CK => Clk, Q => DRAM_DIN(18), QN =>
                           n_1019);
   DATAPATH_IxThird_stxB_FORWARD_out_regx19x : DFF_X1 port map( D => 
                           RF_RD2_DATA(19), CK => Clk, Q => DRAM_DIN(19), QN =>
                           n_1020);
   DATAPATH_IxThird_stxB_FORWARD_out_regx20x : DFF_X1 port map( D => 
                           RF_RD2_DATA(20), CK => Clk, Q => DRAM_DIN(20), QN =>
                           n_1021);
   DATAPATH_IxThird_stxB_FORWARD_out_regx21x : DFF_X1 port map( D => 
                           RF_RD2_DATA(21), CK => Clk, Q => DRAM_DIN(21), QN =>
                           n_1022);
   DATAPATH_IxThird_stxB_FORWARD_out_regx22x : DFF_X1 port map( D => 
                           RF_RD2_DATA(22), CK => Clk, Q => DRAM_DIN(22), QN =>
                           n_1023);
   DATAPATH_IxThird_stxB_FORWARD_out_regx23x : DFF_X1 port map( D => 
                           RF_RD2_DATA(23), CK => Clk, Q => DRAM_DIN(23), QN =>
                           n_1024);
   DATAPATH_IxThird_stxB_FORWARD_out_regx24x : DFF_X1 port map( D => 
                           RF_RD2_DATA(24), CK => Clk, Q => DRAM_DIN(24), QN =>
                           n_1025);
   DATAPATH_IxThird_stxB_FORWARD_out_regx25x : DFF_X1 port map( D => 
                           RF_RD2_DATA(25), CK => Clk, Q => DRAM_DIN(25), QN =>
                           n_1026);
   DATAPATH_IxThird_stxB_FORWARD_out_regx26x : DFF_X1 port map( D => 
                           RF_RD2_DATA(26), CK => Clk, Q => DRAM_DIN(26), QN =>
                           n_1027);
   DATAPATH_IxThird_stxB_FORWARD_out_regx27x : DFF_X1 port map( D => 
                           RF_RD2_DATA(27), CK => Clk, Q => DRAM_DIN(27), QN =>
                           n_1028);
   DATAPATH_IxThird_stxB_FORWARD_out_regx28x : DFF_X1 port map( D => 
                           RF_RD2_DATA(28), CK => Clk, Q => DRAM_DIN(28), QN =>
                           n_1029);
   DATAPATH_IxThird_stxB_FORWARD_out_regx29x : DFF_X1 port map( D => 
                           RF_RD2_DATA(29), CK => Clk, Q => DRAM_DIN(29), QN =>
                           n_1030);
   DATAPATH_IxThird_stxB_FORWARD_out_regx30x : DFF_X1 port map( D => 
                           RF_RD2_DATA(30), CK => Clk, Q => DRAM_DIN(30), QN =>
                           n_1031);
   DATAPATH_IxThird_stxB_FORWARD_out_regx31x : DFF_X1 port map( D => 
                           RF_RD2_DATA(31), CK => Clk, Q => DRAM_DIN(31), QN =>
                           n_1032);
   DATAPATH_IxFourth_stxLMD_out_regx0x : DFF_X1 port map( D => DRAM_DOUT(0), CK
                           => Clk, Q => RF_WR_DATA(0), QN => n_1033);
   DATAPATH_IxFourth_stxLMD_out_regx1x : DFF_X1 port map( D => DRAM_DOUT(1), CK
                           => Clk, Q => RF_WR_DATA(1), QN => n_1034);
   DATAPATH_IxFourth_stxLMD_out_regx2x : DFF_X1 port map( D => DRAM_DOUT(2), CK
                           => Clk, Q => RF_WR_DATA(2), QN => n_1035);
   DATAPATH_IxFourth_stxLMD_out_regx3x : DFF_X1 port map( D => DRAM_DOUT(3), CK
                           => Clk, Q => RF_WR_DATA(3), QN => n_1036);
   DATAPATH_IxFourth_stxLMD_out_regx4x : DFF_X1 port map( D => DRAM_DOUT(4), CK
                           => Clk, Q => RF_WR_DATA(4), QN => n_1037);
   DATAPATH_IxFourth_stxLMD_out_regx5x : DFF_X1 port map( D => DRAM_DOUT(5), CK
                           => Clk, Q => RF_WR_DATA(5), QN => n_1038);
   DATAPATH_IxFourth_stxLMD_out_regx6x : DFF_X1 port map( D => DRAM_DOUT(6), CK
                           => Clk, Q => RF_WR_DATA(6), QN => n_1039);
   DATAPATH_IxFourth_stxLMD_out_regx7x : DFF_X1 port map( D => DRAM_DOUT(7), CK
                           => Clk, Q => RF_WR_DATA(7), QN => n_1040);
   DATAPATH_IxFourth_stxLMD_out_regx8x : DFF_X1 port map( D => DRAM_DOUT(8), CK
                           => Clk, Q => RF_WR_DATA(8), QN => n_1041);
   DATAPATH_IxFourth_stxLMD_out_regx9x : DFF_X1 port map( D => DRAM_DOUT(9), CK
                           => Clk, Q => RF_WR_DATA(9), QN => n_1042);
   DATAPATH_IxFourth_stxLMD_out_regx10x : DFF_X1 port map( D => DRAM_DOUT(10), 
                           CK => Clk, Q => RF_WR_DATA(10), QN => n_1043);
   DATAPATH_IxFourth_stxLMD_out_regx11x : DFF_X1 port map( D => DRAM_DOUT(11), 
                           CK => Clk, Q => RF_WR_DATA(11), QN => n_1044);
   DATAPATH_IxFourth_stxLMD_out_regx12x : DFF_X1 port map( D => DRAM_DOUT(12), 
                           CK => Clk, Q => RF_WR_DATA(12), QN => n_1045);
   DATAPATH_IxFourth_stxLMD_out_regx13x : DFF_X1 port map( D => DRAM_DOUT(13), 
                           CK => Clk, Q => RF_WR_DATA(13), QN => n_1046);
   DATAPATH_IxFourth_stxLMD_out_regx14x : DFF_X1 port map( D => DRAM_DOUT(14), 
                           CK => Clk, Q => RF_WR_DATA(14), QN => n_1047);
   DATAPATH_IxFourth_stxLMD_out_regx15x : DFF_X1 port map( D => DRAM_DOUT(15), 
                           CK => Clk, Q => RF_WR_DATA(15), QN => n_1048);
   DATAPATH_IxFourth_stxLMD_out_regx16x : DFF_X1 port map( D => DRAM_DOUT(16), 
                           CK => Clk, Q => RF_WR_DATA(16), QN => n_1049);
   DATAPATH_IxFourth_stxLMD_out_regx17x : DFF_X1 port map( D => DRAM_DOUT(17), 
                           CK => Clk, Q => RF_WR_DATA(17), QN => n_1050);
   DATAPATH_IxFourth_stxLMD_out_regx18x : DFF_X1 port map( D => DRAM_DOUT(18), 
                           CK => Clk, Q => RF_WR_DATA(18), QN => n_1051);
   DATAPATH_IxFourth_stxLMD_out_regx19x : DFF_X1 port map( D => DRAM_DOUT(19), 
                           CK => Clk, Q => RF_WR_DATA(19), QN => n_1052);
   DATAPATH_IxFourth_stxLMD_out_regx20x : DFF_X1 port map( D => DRAM_DOUT(20), 
                           CK => Clk, Q => RF_WR_DATA(20), QN => n_1053);
   DATAPATH_IxFourth_stxLMD_out_regx21x : DFF_X1 port map( D => DRAM_DOUT(21), 
                           CK => Clk, Q => RF_WR_DATA(21), QN => n_1054);
   DATAPATH_IxFourth_stxLMD_out_regx22x : DFF_X1 port map( D => DRAM_DOUT(22), 
                           CK => Clk, Q => RF_WR_DATA(22), QN => n_1055);
   DATAPATH_IxFourth_stxLMD_out_regx23x : DFF_X1 port map( D => DRAM_DOUT(23), 
                           CK => Clk, Q => RF_WR_DATA(23), QN => n_1056);
   DATAPATH_IxFourth_stxLMD_out_regx24x : DFF_X1 port map( D => DRAM_DOUT(24), 
                           CK => Clk, Q => RF_WR_DATA(24), QN => n_1057);
   DATAPATH_IxFourth_stxLMD_out_regx25x : DFF_X1 port map( D => DRAM_DOUT(25), 
                           CK => Clk, Q => RF_WR_DATA(25), QN => n_1058);
   DATAPATH_IxFourth_stxLMD_out_regx26x : DFF_X1 port map( D => DRAM_DOUT(26), 
                           CK => Clk, Q => RF_WR_DATA(26), QN => n_1059);
   DATAPATH_IxFourth_stxLMD_out_regx27x : DFF_X1 port map( D => DRAM_DOUT(27), 
                           CK => Clk, Q => RF_WR_DATA(27), QN => n_1060);
   DATAPATH_IxFourth_stxLMD_out_regx28x : DFF_X1 port map( D => DRAM_DOUT(28), 
                           CK => Clk, Q => RF_WR_DATA(28), QN => n_1061);
   DATAPATH_IxFourth_stxLMD_out_regx29x : DFF_X1 port map( D => DRAM_DOUT(29), 
                           CK => Clk, Q => RF_WR_DATA(29), QN => n_1062);
   DATAPATH_IxFourth_stxLMD_out_regx30x : DFF_X1 port map( D => DRAM_DOUT(30), 
                           CK => Clk, Q => RF_WR_DATA(30), QN => n_1063);
   DATAPATH_IxFourth_stxLMD_out_regx31x : DFF_X1 port map( D => DRAM_DOUT(31), 
                           CK => Clk, Q => RF_WR_DATA(31), QN => n_1064);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx24x : DFF_X1 port map( D => n696, CK =>
                           Clk, Q => RF_RD2_ADD(4), QN => n717);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx23x : DFF_X1 port map( D => n695, CK =>
                           Clk, Q => RF_RD2_ADD(3), QN => n716);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx22x : DFF_X1 port map( D => n694, CK =>
                           Clk, Q => RF_RD2_ADD(2), QN => n715);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx21x : DFF_X1 port map( D => n693, CK =>
                           Clk, Q => RF_RD2_ADD(1), QN => n714);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx20x : DFF_X1 port map( D => n692, CK =>
                           Clk, Q => RF_RD2_ADD(0), QN => n713);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx19x : DFF_X1 port map( D => n691, CK =>
                           Clk, Q => RF_RD1_ADD(4), QN => n712);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx18x : DFF_X1 port map( D => n690, CK =>
                           Clk, Q => RF_RD1_ADD(3), QN => n711);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx17x : DFF_X1 port map( D => n689, CK =>
                           Clk, Q => RF_RD1_ADD(2), QN => n710);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx16x : DFF_X1 port map( D => n688, CK =>
                           Clk, Q => RF_RD1_ADD(1), QN => n709);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx15x : DFF_X1 port map( D => n687, CK =>
                           Clk, Q => RF_RD1_ADD(0), QN => n708);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx11x : DFF_X1 port map( D => n686, CK =>
                           Clk, Q => DATAPATH_IxINSTR_11_port, QN => n707);
   DATAPATH_IxSecond_stxWRADD_d1_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_11_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, QN => n_1065);
   DATAPATH_IxSecond_stxWRADD_d2_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_4_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_4_port, QN => n_1066);
   DATAPATH_IxSecond_stxWRADD_d3_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_4_port, CK => Clk, Q => 
                           RF_WR_ADD(4), QN => n_1067);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx10x : DFF_X1 port map( D => n685, CK =>
                           Clk, Q => DATAPATH_IxINSTR_10_port, QN => n706);
   DATAPATH_IxSecond_stxWRADD_d1_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_10_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, QN => n_1068);
   DATAPATH_IxSecond_stxWRADD_d2_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_3_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_3_port, QN => n_1069);
   DATAPATH_IxSecond_stxWRADD_d3_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_3_port, CK => Clk, Q => 
                           RF_WR_ADD(3), QN => n_1070);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx9x : DFF_X1 port map( D => n684, CK => 
                           Clk, Q => DATAPATH_IxINSTR_9_port, QN => n705);
   DATAPATH_IxSecond_stxWRADD_d1_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_9_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, QN => n_1071);
   DATAPATH_IxSecond_stxWRADD_d2_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_2_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_2_port, QN => n_1072);
   DATAPATH_IxSecond_stxWRADD_d3_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_2_port, CK => Clk, Q => 
                           RF_WR_ADD(2), QN => n_1073);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx8x : DFF_X1 port map( D => n683, CK => 
                           Clk, Q => DATAPATH_IxINSTR_8_port, QN => n704);
   DATAPATH_IxSecond_stxWRADD_d1_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_8_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, QN => n_1074);
   DATAPATH_IxSecond_stxWRADD_d2_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_1_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_1_port, QN => n_1075);
   DATAPATH_IxSecond_stxWRADD_d3_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_1_port, CK => Clk, Q => 
                           RF_WR_ADD(1), QN => n_1076);
   DATAPATH_IxFirst_stxIR_LATCH_out_regx7x : DFF_X1 port map( D => n682, CK => 
                           Clk, Q => DATAPATH_IxINSTR_7_port, QN => n703);
   DATAPATH_IxSecond_stxWRADD_d1_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxINSTR_7_port, CK => Clk, Q => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, QN => n_1077);
   DATAPATH_IxSecond_stxWRADD_d2_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxSecond_stxWRADD_d1_0_port, CK => Clk, Q 
                           => DATAPATH_IxWR_ADD_MEM_fu_0_port, QN => n_1078);
   DATAPATH_IxSecond_stxWRADD_d3_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxWR_ADD_MEM_fu_0_port, CK => Clk, Q => 
                           RF_WR_ADD(0), QN => n_1079);
   DATAPATH_IxFirst_stxPC_regx2x : DFF_X1 port map( D => n777, CK => Clk, Q => 
                           IRAM_ADD_2_port, QN => n718);
   DATAPATH_IxFirst_stxPC_regx3x : DFF_X1 port map( D => n776, CK => Clk, Q => 
                           IRAM_ADD_3_port, QN => n719);
   DATAPATH_IxFirst_stxPC_regx4x : DFF_X1 port map( D => n775, CK => Clk, Q => 
                           IRAM_ADD_4_port, QN => n720);
   DATAPATH_IxFirst_stxPC_regx5x : DFF_X1 port map( D => n774, CK => Clk, Q => 
                           IRAM_ADD_5_port, QN => n721);
   DATAPATH_IxFirst_stxPC_regx6x : DFF_X1 port map( D => n773, CK => Clk, Q => 
                           IRAM_ADD_6_port, QN => n722);
   DATAPATH_IxFirst_stxPC_regx7x : DFF_X1 port map( D => n772, CK => Clk, Q => 
                           IRAM_ADD_7_port, QN => n723);
   DATAPATH_IxFirst_stxPC_regx8x : DFF_X1 port map( D => n771, CK => Clk, Q => 
                           IRAM_ADD_8_port, QN => n724);
   DATAPATH_IxFirst_stxPC_regx9x : DFF_X1 port map( D => n770, CK => Clk, Q => 
                           IRAM_ADD_9_port, QN => n725);
   DATAPATH_IxFirst_stxPC_regx10x : DFF_X1 port map( D => n769, CK => Clk, Q =>
                           IRAM_ADD_10_port, QN => n726);
   DATAPATH_IxFirst_stxPC_regx11x : DFF_X1 port map( D => n768, CK => Clk, Q =>
                           IRAM_ADD_11_port, QN => n727);
   DATAPATH_IxFirst_stxPC_regx1x : DFF_X1 port map( D => n673, CK => Clk, Q => 
                           DATAPATH_IxPC4_1_port, QN => n668);
   DATAPATH_IxFirst_stxPC_regx0x : DFF_X1 port map( D => n697, CK => Clk, Q => 
                           DATAPATH_IxPC4_0_port, QN => n667);
   DATAPATH_IxFirst_stxPC_regx12x : DFF_X1 port map( D => n767, CK => Clk, Q =>
                           IRAM_ADD_12_port, QN => n728);
   DATAPATH_IxFirst_stxPC_regx13x : DFF_X1 port map( D => n766, CK => Clk, Q =>
                           IRAM_ADD_13_port, QN => n729);
   DATAPATH_IxFirst_stxPC_regx14x : DFF_X1 port map( D => n765, CK => Clk, Q =>
                           IRAM_ADD_14_port, QN => n730);
   DATAPATH_IxFirst_stxPC_regx15x : DFF_X1 port map( D => n764, CK => Clk, Q =>
                           IRAM_ADD_15_port, QN => n731);
   DATAPATH_IxFirst_stxPC_regx16x : DFF_X1 port map( D => n763, CK => Clk, Q =>
                           IRAM_ADD_16_port, QN => n732);
   DATAPATH_IxFirst_stxPC_regx17x : DFF_X1 port map( D => n762, CK => Clk, Q =>
                           IRAM_ADD_17_port, QN => n733);
   DATAPATH_IxFirst_stxPC_regx18x : DFF_X1 port map( D => n761, CK => Clk, Q =>
                           IRAM_ADD_18_port, QN => n734);
   DATAPATH_IxFirst_stxPC_regx19x : DFF_X1 port map( D => n760, CK => Clk, Q =>
                           IRAM_ADD_19_port, QN => n735);
   DATAPATH_IxFirst_stxPC_regx20x : DFF_X1 port map( D => n759, CK => Clk, Q =>
                           IRAM_ADD_20_port, QN => n736);
   DATAPATH_IxFirst_stxPC_regx21x : DFF_X1 port map( D => n758, CK => Clk, Q =>
                           IRAM_ADD_21_port, QN => n737);
   DATAPATH_IxFirst_stxPC_regx22x : DFF_X1 port map( D => n757, CK => Clk, Q =>
                           IRAM_ADD_22_port, QN => n738);
   DATAPATH_IxFirst_stxPC_regx23x : DFF_X1 port map( D => n756, CK => Clk, Q =>
                           IRAM_ADD_23_port, QN => n739);
   DATAPATH_IxFirst_stxPC_regx24x : DFF_X1 port map( D => n755, CK => Clk, Q =>
                           IRAM_ADD_24_port, QN => n740);
   DATAPATH_IxFirst_stxPC_regx25x : DFF_X1 port map( D => n754, CK => Clk, Q =>
                           IRAM_ADD_25_port, QN => n741);
   DATAPATH_IxFirst_stxPC_regx26x : DFF_X1 port map( D => n753, CK => Clk, Q =>
                           IRAM_ADD_26_port, QN => n742);
   DATAPATH_IxFirst_stxPC_regx27x : DFF_X1 port map( D => n752, CK => Clk, Q =>
                           IRAM_ADD_27_port, QN => n743);
   DATAPATH_IxFirst_stxPC_regx28x : DFF_X1 port map( D => n751, CK => Clk, Q =>
                           IRAM_ADD_28_port, QN => n744);
   DATAPATH_IxFirst_stxPC_regx29x : DFF_X1 port map( D => n750, CK => Clk, Q =>
                           IRAM_ADD_29_port, QN => n745);
   DATAPATH_IxFirst_stxPC_regx30x : DFF_X1 port map( D => n749, CK => Clk, Q =>
                           IRAM_ADD_30_port, QN => n746);
   DATAPATH_IxFirst_stxPC_regx31x : DFF_X1 port map( D => n748, CK => Clk, Q =>
                           IRAM_ADD_31_port, QN => n747);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx12x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_12_port, CK => Clk, Q 
                           => DRAM_ADD(12), QN => n_1080);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx16x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_16_port, CK => Clk, Q 
                           => DRAM_ADD(16), QN => n_1081);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx17x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_17_port, CK => Clk, Q 
                           => DRAM_ADD(17), QN => n_1082);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx0x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_0_port, CK => Clk, Q 
                           => DRAM_ADD(0), QN => n_1083);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx10x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_10_port, CK => Clk, Q 
                           => DRAM_ADD(10), QN => n_1084);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx14x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_14_port, CK => Clk, Q 
                           => DRAM_ADD(14), QN => n_1085);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx15x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_15_port, CK => Clk, Q 
                           => DRAM_ADD(15), QN => n_1086);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx31x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_31_port, CK => Clk, Q 
                           => DRAM_ADD(31), QN => n_1087);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx1x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_1_port, CK => Clk, Q 
                           => DRAM_ADD(1), QN => n_1088);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx2x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_2_port, CK => Clk, Q 
                           => DRAM_ADD(2), QN => n_1089);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx3x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_3_port, CK => Clk, Q 
                           => DRAM_ADD(3), QN => n_1090);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx8x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_8_port, CK => Clk, Q 
                           => DRAM_ADD(8), QN => n_1091);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx9x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_9_port, CK => Clk, Q 
                           => DRAM_ADD(9), QN => n_1092);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx28x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_28_port, CK => Clk, Q 
                           => DRAM_ADD(28), QN => n_1093);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx29x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_29_port, CK => Clk, Q 
                           => DRAM_ADD(29), QN => n_1094);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx30x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_30_port, CK => Clk, Q 
                           => DRAM_ADD(30), QN => n_1095);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx4x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_4_port, CK => Clk, Q 
                           => DRAM_ADD(4), QN => n_1096);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx5x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_5_port, CK => Clk, Q 
                           => DRAM_ADD(5), QN => n_1097);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx6x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_6_port, CK => Clk, Q 
                           => DRAM_ADD(6), QN => n_1098);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx7x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_7_port, CK => Clk, Q 
                           => DRAM_ADD(7), QN => n_1099);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx11x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_11_port, CK => Clk, Q 
                           => DRAM_ADD(11), QN => n_1100);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx13x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_13_port, CK => Clk, Q 
                           => DRAM_ADD(13), QN => n_1101);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx18x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_18_port, CK => Clk, Q 
                           => DRAM_ADD(18), QN => n_1102);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx19x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_19_port, CK => Clk, Q 
                           => DRAM_ADD(19), QN => n_1103);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx20x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_20_port, CK => Clk, Q 
                           => DRAM_ADD(20), QN => n_1104);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx21x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_21_port, CK => Clk, Q 
                           => DRAM_ADD(21), QN => n_1105);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx22x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_22_port, CK => Clk, Q 
                           => DRAM_ADD(22), QN => n_1106);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx23x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_23_port, CK => Clk, Q 
                           => DRAM_ADD(23), QN => n_1107);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx24x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_24_port, CK => Clk, Q 
                           => DRAM_ADD(24), QN => n_1108);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx25x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_25_port, CK => Clk, Q 
                           => DRAM_ADD(25), QN => n_1109);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx26x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_26_port, CK => Clk, Q 
                           => DRAM_ADD(26), QN => n_1110);
   DATAPATH_IxThird_stxALU_OUT_MEM_regx27x : DFF_X1 port map( D => 
                           DATAPATH_IxThird_stxALU_out_i_27_port, CK => Clk, Q 
                           => DRAM_ADD(27), QN => n_1111);
   U8 : NAND3_X1 port map( A1 => n23, A2 => n24, A3 => n824, ZN => n679);
   U17 : NAND3_X1 port map( A1 => n33, A2 => n24, A3 => n37, ZN => n681);
   U22 : NAND3_X1 port map( A1 => n36, A2 => n853, A3 => IRAM_DOUT(14), ZN => 
                           n24);
   U65 : NAND3_X1 port map( A1 => n65, A2 => n803, A3 => n746, ZN => n70);
   U71 : NAND3_X1 port map( A1 => n72, A2 => n804, A3 => n745, ZN => n74);
   U80 : NAND3_X1 port map( A1 => n79, A2 => n804, A3 => n743, ZN => n82);
   U90 : NAND3_X1 port map( A1 => n87, A2 => n804, A3 => n741, ZN => n91);
   U100 : NAND3_X1 port map( A1 => n95, A2 => n804, A3 => n739, ZN => n99);
   U112 : NAND3_X1 port map( A1 => IRAM_ADD_20_port, A2 => IRAM_ADD_19_port, A3
                           => n109, ZN => n100);
   U119 : NAND3_X1 port map( A1 => n109, A2 => n804, A3 => n735, ZN => n114);
   U129 : NAND3_X1 port map( A1 => n118, A2 => n804, A3 => n733, ZN => n122);
   U139 : NAND3_X1 port map( A1 => n126, A2 => n804, A3 => n731, ZN => n130);
   U149 : NAND3_X1 port map( A1 => n134, A2 => n804, A3 => n729, ZN => n138);
   U159 : NAND3_X1 port map( A1 => n142, A2 => n804, A3 => n727, ZN => n146);
   U169 : NAND3_X1 port map( A1 => n150, A2 => n804, A3 => n725, ZN => n154);
   U179 : NAND3_X1 port map( A1 => n158, A2 => n804, A3 => n723, ZN => n162);
   U189 : NAND3_X1 port map( A1 => n166, A2 => n804, A3 => n721, ZN => n170);
   U199 : NAND3_X1 port map( A1 => n803, A2 => IRAM_ADD_2_port, A3 => n719, ZN 
                           => n177);
   U213 : XOR2_X1 port map( A => n186, B => n187, Z => n184);
   U215 : NAND3_X1 port map( A1 => n795, A2 => n936, A3 => RF_RD1_DATA(9), ZN 
                           => n181);
   U221 : XOR2_X1 port map( A => n191, B => n881, Z => n200);
   U222 : NAND3_X1 port map( A1 => n796, A2 => n937, A3 => RF_RD1_DATA(8), ZN 
                           => n198);
   U230 : XOR2_X1 port map( A => n216, B => n217, Z => n214);
   U232 : XOR2_X1 port map( A => n221, B => n217, Z => n213);
   U240 : XOR2_X1 port map( A => n219, B => n232, Z => n231);
   U242 : XOR2_X1 port map( A => n222, B => n232, Z => n230);
   U250 : NAND3_X1 port map( A1 => n796, A2 => n814, A3 => RF_RD1_DATA(5), ZN 
                           => n239);
   U256 : XOR2_X1 port map( A => n215, B => n252, Z => n251);
   U257 : NAND3_X1 port map( A1 => n796, A2 => n815, A3 => RF_RD1_DATA(4), ZN 
                           => n249);
   U265 : XOR2_X1 port map( A => n263, B => n264, Z => n261);
   U267 : XOR2_X1 port map( A => n263, B => n268, Z => n259);
   U272 : NAND3_X1 port map( A1 => n796, A2 => n925, A3 => n781, ZN => n274);
   U280 : XOR2_X1 port map( A => n287, B => n288, Z => n285);
   U281 : XOR2_X1 port map( A => n289, B => n287, Z => n283);
   U287 : XOR2_X1 port map( A => n266, B => n297, Z => n296);
   U289 : XOR2_X1 port map( A => n269, B => n297, Z => n295);
   U293 : XOR2_X1 port map( A => n307, B => n308, Z => n306);
   U296 : NAND3_X1 port map( A1 => n796, A2 => n926, A3 => RF_RD1_DATA(29), ZN 
                           => n304);
   U301 : XOR2_X1 port map( A => n286, B => n319, Z => n318);
   U312 : XOR2_X1 port map( A => n329, B => n330, Z => n327);
   U314 : XOR2_X1 port map( A => n334, B => n329, Z => n325);
   U322 : XOR2_X1 port map( A => n331, B => n343, Z => n342);
   U324 : XOR2_X1 port map( A => n343, B => n335, Z => n341);
   U333 : NAND3_X1 port map( A1 => n795, A2 => n928, A3 => RF_RD1_DATA(25), ZN 
                           => n352);
   U339 : XOR2_X1 port map( A => n326, B => n366, Z => n365);
   U348 : XOR2_X1 port map( A => n376, B => n377, Z => n375);
   U350 : XOR2_X1 port map( A => n381, B => n377, Z => n372);
   U358 : XOR2_X1 port map( A => n379, B => n392, Z => n391);
   U360 : NAND3_X1 port map( A1 => n395, A2 => n890, A3 => n893, ZN => n394);
   U361 : XOR2_X1 port map( A => n382, B => n392, Z => n390);
   U370 : NAND3_X1 port map( A1 => n795, A2 => n930, A3 => RF_RD1_DATA(21), ZN 
                           => n402);
   U376 : XOR2_X1 port map( A => n373, B => n416, Z => n415);
   U386 : XOR2_X1 port map( A => n424, B => n298, Z => n423);
   U395 : XOR2_X1 port map( A => n437, B => n875, Z => n435);
   U397 : XOR2_X1 port map( A => n875, B => n442, Z => n433);
   U404 : XOR2_X1 port map( A => n871, B => n874, Z => n450);
   U407 : XOR2_X1 port map( A => n871, B => n873, Z => n449);
   U417 : NAND3_X1 port map( A1 => n796, A2 => n932, A3 => RF_RD1_DATA(17), ZN 
                           => n462);
   U423 : XOR2_X1 port map( A => n436, B => n476, Z => n475);
   U432 : XOR2_X1 port map( A => n486, B => n487, Z => n485);
   U434 : XOR2_X1 port map( A => n491, B => n487, Z => n482);
   U442 : XOR2_X1 port map( A => n489, B => n502, Z => n501);
   U444 : XOR2_X1 port map( A => n492, B => n502, Z => n500);
   U452 : NAND3_X1 port map( A1 => n795, A2 => n934, A3 => RF_RD1_DATA(13), ZN 
                           => n509);
   U458 : XOR2_X1 port map( A => n483, B => n523, Z => n522);
   U470 : XOR2_X1 port map( A => n532, B => n533, Z => n531);
   U472 : XOR2_X1 port map( A => n532, B => n537, Z => n529);
   U479 : XOR2_X1 port map( A => n534, B => n546, Z => n545);
   U483 : XOR2_X1 port map( A => n538, B => n546, Z => n544);
   U489 : NAND3_X1 port map( A1 => n702, A2 => n945, A3 => n701, ZN => n558);
   U490 : XOR2_X1 port map( A => n560, B => n262, Z => n555);
   U500 : XOR2_X1 port map( A => n566, B => n567, Z => n565);
   U501 : XOR2_X1 port map( A => n568, B => n276, Z => n567);
   U511 : XOR2_X1 port map( A => n311, B => n310, Z => n319);
   U531 : XOR2_X1 port map( A => n784, B => n926, Z => n582);
   U562 : XOR2_X1 port map( A => n467, B => n468, Z => n476);
   U617 : XOR2_X1 port map( A => n426, B => n425, Z => n560);
   U620 : XOR2_X1 port map( A => n270, B => n271, Z => n297);
   U621 : XOR2_X1 port map( A => n784, B => n818, Z => n271);
   U624 : XOR2_X1 port map( A => n784, B => n816, Z => n638);
   U625 : XOR2_X1 port map( A => n786, B => RF_RD1_DATA(3), Z => n637);
   U626 : XOR2_X1 port map( A => n244, B => n245, Z => n252);
   U627 : XOR2_X1 port map( A => n784, B => n815, Z => n245);
   U629 : XOR2_X1 port map( A => n787, B => n920, Z => n244);
   U631 : XOR2_X1 port map( A => n224, B => n223, Z => n232);
   U632 : XOR2_X1 port map( A => n784, B => RF_RD2_DATA(6), Z => n223);
   U635 : XOR2_X1 port map( A => n784, B => RF_RD2_DATA(7), Z => n629);
   U636 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(7), Z => n628);
   U640 : XOR2_X1 port map( A => n787, B => n916, Z => n189);
   U642 : XOR2_X1 port map( A => n784, B => n937, Z => n188);
   U650 : XOR2_X1 port map( A => n784, B => RF_RD2_DATA(10), Z => n648);
   U651 : XOR2_X1 port map( A => n784, B => RF_RD2_DATA(11), Z => n621);
   U652 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(11), Z => n620);
   U653 : XOR2_X1 port map( A => n515, B => n514, Z => n523);
   U654 : XOR2_X1 port map( A => n784, B => n935, Z => n514);
   U656 : XOR2_X1 port map( A => n787, B => n912, Z => n515);
   U658 : XOR2_X1 port map( A => n494, B => n493, Z => n502);
   U659 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(14), Z => n493);
   U662 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(15), Z => n612);
   U663 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(15), Z => n611);
   U666 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(19), Z => n606);
   U667 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(19), Z => n607);
   U672 : XOR2_X1 port map( A => n787, B => n908, Z => n467);
   U674 : XOR2_X1 port map( A => n783, B => n933, Z => n468);
   U683 : XOR2_X1 port map( A => n787, B => n906, Z => n651);
   U686 : XOR2_X1 port map( A => n893, B => n395, Z => n416);
   U687 : XOR2_X1 port map( A => n787, B => n904, Z => n395);
   U690 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(20), Z => n407);
   U691 : XOR2_X1 port map( A => n384, B => n383, Z => n392);
   U692 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(22), Z => n383);
   U695 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(23), Z => n598);
   U696 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(23), Z => n597);
   U697 : XOR2_X1 port map( A => n358, B => n357, Z => n366);
   U698 : XOR2_X1 port map( A => n783, B => n929, Z => n357);
   U700 : XOR2_X1 port map( A => n787, B => n900, Z => n358);
   U706 : XOR2_X1 port map( A => n787, B => RF_RD1_DATA(26), Z => n654);
   U707 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(26), Z => n655);
   U708 : XOR2_X1 port map( A => n783, B => RF_RD2_DATA(27), Z => n592);
   U710 : XOR2_X1 port map( A => n786, B => RF_RD1_DATA(27), Z => n591);
   U730 : NAND3_X1 port map( A1 => IRAM_DOUT(1), A2 => IRAM_DOUT(0), A3 => 
                           IRAM_DOUT(5), ZN => n663);
   RF_WR_EN <= '0';
   DRAM_RE <= '0';
   DRAM_WE <= '0';
   RF_RD1_EN <= '0';
   RF_RD2_EN <= '0';
   U209 : AOI21_X2 port map( B1 => n939, B2 => n698, A => n840, ZN => n83);
   CU_Ixstate_var_regx1x : DFFR_X1 port map( D => CU_IxN53, CK => Clk, RN => 
                           Rst, Q => n939, QN => n_1112);
   CU_IxaluOpcode3_regx3x : DFF_X1 port map( D => n674, CK => Clk, Q => n947, 
                           QN => n702);
   CU_IxaluOpcode3_regx2x : DFF_X1 port map( D => n675, CK => Clk, Q => n_1113,
                           QN => n701);
   CU_IxaluOpcode3_regx1x : DFF_X1 port map( D => n676, CK => Clk, Q => n945, 
                           QN => n700);
   CU_IxaluOpcode3_regx0x : DFF_X1 port map( D => n677, CK => Clk, Q => n944, 
                           QN => n699);
   CU_IxaluOpcode2_regx1x : DFF_X1 port map( D => n680, CK => Clk, Q => n_1114,
                           QN => n671);
   CU_IxaluOpcode2_regx2x : DFF_X1 port map( D => n679, CK => Clk, Q => n_1115,
                           QN => n670);
   CU_IxaluOpcode2_regx0x : DFF_X1 port map( D => n681, CK => Clk, Q => n940, 
                           QN => n672);
   CU_IxaluOpcode2_regx3x : DFF_X1 port map( D => n678, CK => Clk, Q => n_1116,
                           QN => n669);
   U742 : OAI21_X2 port map( B1 => n556, B2 => n946, A => n558, ZN => n204);
   U743 : BUF_X1 port map( A => RF_RD2_DATA(1), Z => n820);
   U744 : BUF_X1 port map( A => RF_RD2_DATA(0), Z => n822);
   U745 : INV_X1 port map( A => n550, ZN => n880);
   U746 : INV_X1 port map( A => n610, ZN => n871);
   U747 : INV_X1 port map( A => n236, ZN => n883);
   U748 : INV_X1 port map( A => n504, ZN => n877);
   U749 : INV_X1 port map( A => n812, ZN => n803);
   U750 : INV_X1 port map( A => n812, ZN => n804);
   U751 : XNOR2_X1 port map( A => n242, B => n243, ZN => n241);
   U752 : AOI21_X1 port map( B1 => n236, B2 => n884, A => n233, ZN => n242);
   U753 : XNOR2_X1 port map( A => n885, B => n424, ZN => n422);
   U754 : XNOR2_X1 port map( A => n512, B => n513, ZN => n511);
   U755 : AOI21_X1 port map( B1 => n504, B2 => n878, A => n506, ZN => n512);
   U756 : INV_X1 port map( A => n345, ZN => n868);
   U757 : BUF_X1 port map( A => n585, Z => n786);
   U758 : BUF_X1 port map( A => n585, Z => n785);
   U759 : BUF_X1 port map( A => n585, Z => n787);
   U760 : OAI22_X1 port map( A1 => n286, A2 => n569, B1 => n866, B2 => n570, ZN
                           => n276);
   U761 : XNOR2_X1 port map( A => n573, B => n572, ZN => n569);
   U762 : XNOR2_X1 port map( A => n571, B => n572, ZN => n570);
   U763 : NOR2_X1 port map( A1 => n271, A2 => n270, ZN => n267);
   U764 : NOR2_X1 port map( A1 => n536, A2 => n879, ZN => n546);
   U765 : INV_X1 port map( A => n535, ZN => n879);
   U766 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(5), ZN => n635);
   U767 : AOI22_X1 port map( A1 => n415, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN287, B2 => n798, ZN => 
                           n414);
   U768 : AOI22_X1 port map( A1 => n318, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN295, B2 => n798, ZN => 
                           n317);
   U769 : NAND2_X1 port map( A1 => n188, A2 => n189, ZN => n550);
   U770 : BUF_X1 port map( A => n586, Z => n783);
   U771 : BUF_X1 port map( A => n586, Z => n782);
   U772 : NOR2_X1 port map( A1 => n872, A2 => n439, ZN => n610);
   U773 : BUF_X1 port map( A => n586, Z => n784);
   U774 : NAND2_X1 port map( A1 => n468, A2 => n467, ZN => n457);
   U775 : NAND2_X1 port map( A1 => n245, A2 => n244, ZN => n236);
   U776 : NAND2_X1 port map( A1 => n515, A2 => n514, ZN => n504);
   U777 : INV_X1 port map( A => n373, ZN => n870);
   U778 : INV_X1 port map( A => n262, ZN => n892);
   U779 : XNOR2_X1 port map( A => n465, B => n466, ZN => n464);
   U780 : AOI21_X1 port map( B1 => n457, B2 => n876, A => n453, ZN => n465);
   U781 : INV_X1 port map( A => n286, ZN => n866);
   U782 : XNOR2_X1 port map( A => n355, B => n356, ZN => n354);
   U783 : AOI21_X1 port map( B1 => n345, B2 => n869, A => n347, ZN => n355);
   U784 : INV_X1 port map( A => n326, ZN => n869);
   U785 : INV_X1 port map( A => n436, ZN => n876);
   U786 : NAND2_X1 port map( A1 => n300, A2 => n886, ZN => n424);
   U787 : INV_X1 port map( A => n299, ZN => n886);
   U788 : NOR2_X1 port map( A1 => n466, A2 => n871, ZN => n609);
   U789 : NAND2_X1 port map( A1 => n887, A2 => n235, ZN => n243);
   U790 : INV_X1 port map( A => n234, ZN => n887);
   U791 : NAND2_X1 port map( A1 => n889, A2 => n505, ZN => n513);
   U792 : INV_X1 port map( A => n503, ZN => n889);
   U793 : INV_X1 port map( A => n605, ZN => n875);
   U794 : NAND2_X1 port map( A1 => n888, A2 => n549, ZN => n186);
   U795 : INV_X1 port map( A => n547, ZN => n888);
   U796 : INV_X1 port map( A => n645, ZN => n881);
   U797 : OAI21_X1 port map( B1 => n188, B2 => n189, A => n550, ZN => n645);
   U798 : INV_X1 port map( A => n301, ZN => n885);
   U799 : INV_X1 port map( A => n441, ZN => n872);
   U800 : XNOR2_X1 port map( A => n575, B => n574, ZN => n572);
   U801 : AOI21_X1 port map( B1 => n289, B2 => n583, A => n891, ZN => n573);
   U802 : AOI21_X1 port map( B1 => n288, B2 => n583, A => n891, ZN => n571);
   U803 : OAI22_X1 port map( A1 => n188, A2 => n189, B1 => n880, B2 => n191, ZN
                           => n187);
   U804 : OAI21_X1 port map( B1 => n378, B2 => n379, A => n380, ZN => n376);
   U805 : OAI21_X1 port map( B1 => n492, B2 => n488, A => n490, ZN => n491);
   U806 : AOI21_X1 port map( B1 => n332, B2 => n335, A => n333, ZN => n334);
   U807 : OAI21_X1 port map( B1 => n873, B2 => n439, A => n441, ZN => n442);
   U808 : AOI21_X1 port map( B1 => n265, B2 => n269, A => n267, ZN => n268);
   U809 : AOI21_X1 port map( B1 => n538, B2 => n535, A => n536, ZN => n537);
   U810 : OAI21_X1 port map( B1 => n218, B2 => n219, A => n220, ZN => n216);
   U811 : OAI21_X1 port map( B1 => n439, B2 => n874, A => n441, ZN => n437);
   U812 : AOI21_X1 port map( B1 => n331, B2 => n332, A => n333, ZN => n330);
   U813 : AOI21_X1 port map( B1 => n534, B2 => n535, A => n536, ZN => n533);
   U814 : NOR2_X1 port map( A1 => n333, A2 => n867, ZN => n343);
   U815 : INV_X1 port map( A => n332, ZN => n867);
   U816 : OAI21_X1 port map( B1 => n347, B2 => n344, A => n346, ZN => n335);
   U817 : OAI21_X1 port map( B1 => n298, B2 => n299, A => n300, ZN => n266);
   U818 : OAI21_X1 port map( B1 => n299, B2 => n301, A => n300, ZN => n269);
   U819 : OAI21_X1 port map( B1 => n234, B2 => n236, A => n235, ZN => n222);
   U820 : OAI21_X1 port map( B1 => n503, B2 => n504, A => n505, ZN => n489);
   U821 : OAI21_X1 port map( B1 => n398, B2 => n399, A => n393, ZN => n382);
   U822 : NOR2_X1 port map( A1 => n893, A2 => n395, ZN => n398);
   U823 : OAI21_X1 port map( B1 => n547, B2 => n550, A => n549, ZN => n538);
   U824 : OAI21_X1 port map( B1 => n233, B2 => n234, A => n235, ZN => n219);
   U825 : OAI21_X1 port map( B1 => n344, B2 => n345, A => n346, ZN => n331);
   U826 : NOR2_X1 port map( A1 => n467, A2 => n468, ZN => n453);
   U827 : NOR2_X1 port map( A1 => n244, A2 => n245, ZN => n233);
   U828 : OAI21_X1 port map( B1 => n547, B2 => n548, A => n549, ZN => n534);
   U829 : NOR2_X1 port map( A1 => n188, A2 => n189, ZN => n548);
   U830 : OAI21_X1 port map( B1 => n506, B2 => n503, A => n505, ZN => n492);
   U831 : NOR2_X1 port map( A1 => n357, A2 => n358, ZN => n347);
   U832 : NOR2_X1 port map( A1 => n514, A2 => n515, ZN => n506);
   U833 : NAND2_X1 port map( A1 => n358, A2 => n357, ZN => n345);
   U834 : AOI21_X1 port map( B1 => n265, B2 => n266, A => n267, ZN => n264);
   U835 : INV_X1 port map( A => n456, ZN => n873);
   U836 : OAI21_X1 port map( B1 => n454, B2 => n457, A => n455, ZN => n456);
   U837 : NAND2_X1 port map( A1 => n780, A2 => n786, ZN => n575);
   U838 : INV_X1 port map( A => n483, ZN => n878);
   U839 : INV_X1 port map( A => n215, ZN => n884);
   U840 : INV_X1 port map( A => n191, ZN => n882);
   U841 : OAI21_X1 port map( B1 => n488, B2 => n489, A => n490, ZN => n486);
   U842 : OAI21_X1 port map( B1 => n378, B2 => n382, A => n380, ZN => n381);
   U843 : OAI21_X1 port map( B1 => n218, B2 => n222, A => n220, ZN => n221);
   U844 : NAND2_X1 port map( A1 => n393, A2 => n394, ZN => n379);
   U845 : BUF_X1 port map( A => n802, Z => n812);
   U846 : NAND2_X1 port map( A1 => n270, A2 => n271, ZN => n265);
   U847 : BUF_X1 port map( A => n800, Z => n806);
   U848 : BUF_X1 port map( A => n800, Z => n805);
   U849 : BUF_X1 port map( A => n800, Z => n807);
   U850 : INV_X1 port map( A => n584, ZN => n891);
   U851 : BUF_X1 port map( A => n801, Z => n810);
   U852 : BUF_X1 port map( A => n801, Z => n809);
   U853 : BUF_X1 port map( A => n801, Z => n808);
   U854 : BUF_X1 port map( A => n802, Z => n811);
   U855 : NAND2_X1 port map( A1 => n393, A2 => n890, ZN => n405);
   U856 : AND2_X1 port map( A1 => n583, A2 => n584, ZN => n287);
   U857 : INV_X1 port map( A => n452, ZN => n874);
   U858 : OAI21_X1 port map( B1 => n453, B2 => n454, A => n455, ZN => n452);
   U859 : INV_X1 port map( A => n399, ZN => n890);
   U860 : INV_X1 port map( A => n795, ZN => n788);
   U861 : INV_X1 port map( A => n795, ZN => n789);
   U862 : BUF_X1 port map( A => n781, Z => n779);
   U863 : BUF_X1 port map( A => RF_RD1_DATA(31), Z => n780);
   U864 : BUF_X1 port map( A => RF_RD1_DATA(31), Z => n781);
   U865 : OAI22_X1 port map( A1 => n628, A2 => n629, B1 => n630, B2 => n217, ZN
                           => n191);
   U866 : AOI21_X1 port map( B1 => n232, B2 => n631, A => n218, ZN => n630);
   U867 : OAI21_X1 port map( B1 => n632, B2 => n243, A => n235, ZN => n631);
   U868 : AOI21_X1 port map( B1 => n252, B2 => n215, A => n883, ZN => n632);
   U869 : OAI22_X1 port map( A1 => n591, A2 => n592, B1 => n593, B2 => n329, ZN
                           => n286);
   U870 : AOI21_X1 port map( B1 => n343, B2 => n594, A => n333, ZN => n593);
   U871 : OAI21_X1 port map( B1 => n595, B2 => n356, A => n346, ZN => n594);
   U872 : AOI21_X1 port map( B1 => n366, B2 => n326, A => n868, ZN => n595);
   U873 : OAI21_X1 port map( B1 => n656, B2 => n813, A => n946, ZN => n262);
   U874 : OAI22_X1 port map( A1 => n597, A2 => n598, B1 => n599, B2 => n377, ZN
                           => n326);
   U875 : AOI21_X1 port map( B1 => n392, B2 => n600, A => n378, ZN => n599);
   U876 : OAI21_X1 port map( B1 => n601, B2 => n405, A => n393, ZN => n600);
   U877 : AOI22_X1 port map( A1 => n416, A2 => n373, B1 => n893, B2 => n395, ZN
                           => n601);
   U878 : OAI22_X1 port map( A1 => n620, A2 => n621, B1 => n622, B2 => n532, ZN
                           => n483);
   U879 : AOI21_X1 port map( B1 => n546, B2 => n623, A => n536, ZN => n622);
   U880 : OAI21_X1 port map( B1 => n624, B2 => n186, A => n549, ZN => n623);
   U881 : AOI21_X1 port map( B1 => n881, B2 => n191, A => n880, ZN => n624);
   U882 : OAI22_X1 port map( A1 => n637, A2 => n638, B1 => n639, B2 => n263, ZN
                           => n215);
   U883 : AOI21_X1 port map( B1 => n297, B2 => n640, A => n267, ZN => n639);
   U884 : OAI21_X1 port map( B1 => n641, B2 => n424, A => n300, ZN => n640);
   U885 : AOI21_X1 port map( B1 => n560, B2 => n262, A => n885, ZN => n641);
   U886 : OAI22_X1 port map( A1 => n611, A2 => n612, B1 => n613, B2 => n487, ZN
                           => n436);
   U887 : AOI21_X1 port map( B1 => n502, B2 => n614, A => n488, ZN => n613);
   U888 : OAI21_X1 port map( B1 => n615, B2 => n513, A => n505, ZN => n614);
   U889 : AOI21_X1 port map( B1 => n523, B2 => n483, A => n877, ZN => n615);
   U890 : NOR2_X1 port map( A1 => n648, A2 => n647, ZN => n536);
   U891 : XNOR2_X1 port map( A => n458, B => n459, ZN => n466);
   U892 : XNOR2_X1 port map( A => n785, B => n910, ZN => n494);
   U893 : XNOR2_X1 port map( A => n785, B => n918, ZN => n224);
   U894 : XNOR2_X1 port map( A => n785, B => n922, ZN => n270);
   U895 : XNOR2_X1 port map( A => n783, B => n822, ZN => n425);
   U896 : NOR2_X1 port map( A1 => n651, A2 => n652, ZN => n439);
   U897 : NOR2_X1 port map( A1 => n635, A2 => n634, ZN => n234);
   U898 : NOR2_X1 port map( A1 => n618, A2 => n617, ZN => n503);
   U899 : NOR2_X1 port map( A1 => n643, A2 => n644, ZN => n299);
   U900 : NOR2_X1 port map( A1 => n494, A2 => n493, ZN => n488);
   U901 : XNOR2_X1 port map( A => n611, B => n612, ZN => n487);
   U902 : XNOR2_X1 port map( A => n628, B => n629, ZN => n217);
   U903 : NOR2_X1 port map( A1 => n627, A2 => n626, ZN => n547);
   U904 : NOR2_X1 port map( A1 => n224, A2 => n223, ZN => n218);
   U905 : XNOR2_X1 port map( A => n637, B => n638, ZN => n263);
   U906 : XNOR2_X1 port map( A => n620, B => n621, ZN => n532);
   U907 : AOI22_X1 port map( A1 => n309, A2 => n286, B1 => n310, B2 => n311, ZN
                           => n308);
   U908 : OR2_X1 port map( A1 => n311, A2 => n310, ZN => n309);
   U909 : XNOR2_X1 port map( A => n782, B => n820, ZN => n643);
   U910 : OAI22_X1 port map( A1 => n574, A2 => n575, B1 => n576, B2 => n572, ZN
                           => n568);
   U911 : AOI21_X1 port map( B1 => n287, B2 => n577, A => n891, ZN => n576);
   U912 : OAI21_X1 port map( B1 => n579, B2 => n307, A => n580, ZN => n577);
   U913 : AOI22_X1 port map( A1 => n319, A2 => n286, B1 => n310, B2 => n311, ZN
                           => n579);
   U914 : XNOR2_X1 port map( A => n785, B => n914, ZN => n647);
   U915 : XNOR2_X1 port map( A => n607, B => n606, ZN => n605);
   U916 : XNOR2_X1 port map( A => n405, B => n406, ZN => n404);
   U917 : AOI21_X1 port map( B1 => n870, B2 => n407, A => n408, ZN => n406);
   U918 : AOI21_X1 port map( B1 => n893, B2 => n373, A => n395, ZN => n408);
   U919 : OAI221_X1 port map( B1 => n604, B2 => n605, C1 => n606, C2 => n607, A
                           => n608, ZN => n373);
   U920 : AOI21_X1 port map( B1 => n610, B2 => n649, A => n872, ZN => n604);
   U921 : NAND4_X1 port map( A1 => n875, A2 => n436, A3 => n476, A4 => n609, ZN
                           => n608);
   U922 : OAI21_X1 port map( B1 => n466, B2 => n457, A => n455, ZN => n649);
   U923 : NAND2_X1 port map( A1 => n634, A2 => n635, ZN => n235);
   U924 : NAND2_X1 port map( A1 => n617, A2 => n618, ZN => n505);
   U925 : NAND2_X1 port map( A1 => n626, A2 => n627, ZN => n549);
   U926 : NAND2_X1 port map( A1 => n644, A2 => n643, ZN => n300);
   U927 : INV_X1 port map( A => n564, ZN => n946);
   U928 : NAND2_X1 port map( A1 => n652, A2 => n651, ZN => n441);
   U929 : NAND2_X1 port map( A1 => n656, A2 => n262, ZN => n586);
   U930 : NAND2_X1 port map( A1 => n459, A2 => n458, ZN => n455);
   U931 : NAND2_X1 port map( A1 => n647, A2 => n648, ZN => n535);
   U932 : OAI211_X1 port map( C1 => n272, C2 => n925, A => n274, B => n275, ZN 
                           => DATAPATH_IxThird_stxALU_out_i_31_port);
   U933 : AOI221_X1 port map( B1 => n792, B2 => n813, C1 => n780, C2 => n942, A
                           => n941, ZN => n272);
   U934 : AOI22_X1 port map( A1 => n943, A2 => n276, B1 => n781, B2 => n799, ZN
                           => n275);
   U935 : NAND2_X1 port map( A1 => n425, A2 => n426, ZN => n301);
   U936 : NAND4_X1 port map( A1 => n551, A2 => n552, A3 => n553, A4 => n554, ZN
                           => DATAPATH_IxThird_stxALU_out_i_0_port);
   U937 : NAND2_X1 port map( A1 => n822, A2 => n561, ZN => n553);
   U938 : OR3_X1 port map( A1 => n789, A2 => n822, A3 => n924, ZN => n551);
   U939 : AOI22_X1 port map( A1 => DATAPATH_IxThird_stxALU1xN267, A2 => n797, 
                           B1 => n555, B2 => n943, ZN => n554);
   U940 : OR2_X1 port map( A1 => n656, A2 => n892, ZN => n585);
   U941 : INV_X1 port map( A => n83, ZN => n839);
   U942 : NOR2_X1 port map( A1 => n655, A2 => n654, ZN => n333);
   U943 : AOI21_X1 port map( B1 => n948, B2 => n803, A => n83, ZN => n81);
   U944 : AOI21_X1 port map( B1 => n949, B2 => n804, A => n83, ZN => n90);
   U945 : AOI21_X1 port map( B1 => n950, B2 => n804, A => n83, ZN => n98);
   U946 : AOI21_X1 port map( B1 => n951, B2 => n803, A => n83, ZN => n121);
   U947 : AOI21_X1 port map( B1 => n952, B2 => n803, A => n83, ZN => n129);
   U948 : AOI21_X1 port map( B1 => n953, B2 => n803, A => n83, ZN => n137);
   U949 : AOI21_X1 port map( B1 => n954, B2 => n804, A => n83, ZN => n145);
   U950 : AOI21_X1 port map( B1 => n955, B2 => n803, A => n83, ZN => n153);
   U951 : AOI21_X1 port map( B1 => n956, B2 => n803, A => n83, ZN => n161);
   U952 : AOI21_X1 port map( B1 => n957, B2 => n804, A => n83, ZN => n169);
   U953 : XNOR2_X1 port map( A => n785, B => n902, ZN => n384);
   U954 : XNOR2_X1 port map( A => n597, B => n598, ZN => n377);
   U955 : XNOR2_X1 port map( A => n591, B => n592, ZN => n329);
   U956 : NOR2_X1 port map( A1 => n384, A2 => n383, ZN => n378);
   U957 : XNOR2_X1 port map( A => n348, B => n349, ZN => n356);
   U958 : XNOR2_X1 port map( A => n782, B => n925, ZN => n574);
   U959 : OAI21_X1 port map( B1 => n65, B2 => n807, A => n839, ZN => n68);
   U960 : OAI21_X1 port map( B1 => n109, B2 => n806, A => n839, ZN => n112);
   U961 : XNOR2_X1 port map( A => n581, B => n582, ZN => n307);
   U962 : OAI21_X1 port map( B1 => n811, B2 => IRAM_ADD_27_port, A => n81, ZN 
                           => n76);
   U963 : OAI211_X1 port map( C1 => n290, C2 => n204, A => n291, B => n292, ZN 
                           => DATAPATH_IxThird_stxALU_out_i_2_port);
   U964 : OR3_X1 port map( A1 => n788, A2 => n818, A3 => n922, ZN => n291);
   U965 : AOI22_X1 port map( A1 => n818, A2 => n293, B1 => 
                           DATAPATH_IxThird_stxALU1xN269, B2 => n798, ZN => 
                           n292);
   U966 : AOI22_X1 port map( A1 => n295, A2 => n892, B1 => n296, B2 => n262, ZN
                           => n290);
   U967 : OAI211_X1 port map( C1 => n254, C2 => n204, A => n255, B => n256, ZN 
                           => DATAPATH_IxThird_stxALU_out_i_3_port);
   U968 : OR3_X1 port map( A1 => n789, A2 => n816, A3 => n921, ZN => n255);
   U969 : AOI22_X1 port map( A1 => n816, A2 => n257, B1 => 
                           DATAPATH_IxThird_stxALU1xN270, B2 => n799, ZN => 
                           n256);
   U970 : AOI22_X1 port map( A1 => n259, A2 => n892, B1 => n261, B2 => n262, ZN
                           => n254);
   U971 : OAI211_X1 port map( C1 => n417, C2 => n204, A => n418, B => n419, ZN 
                           => DATAPATH_IxThird_stxALU_out_i_1_port);
   U972 : OR3_X1 port map( A1 => n788, A2 => n820, A3 => n923, ZN => n418);
   U973 : AOI22_X1 port map( A1 => n820, A2 => n420, B1 => 
                           DATAPATH_IxThird_stxALU1xN268, B2 => n797, ZN => 
                           n419);
   U974 : AOI22_X1 port map( A1 => n892, A2 => n422, B1 => n423, B2 => n262, ZN
                           => n417);
   U975 : NOR2_X1 port map( A1 => n348, A2 => n349, ZN => n344);
   U976 : NOR2_X1 port map( A1 => n458, A2 => n459, ZN => n454);
   U977 : NOR2_X1 port map( A1 => n602, A2 => n603, ZN => n399);
   U978 : NAND2_X1 port map( A1 => n581, A2 => n582, ZN => n580);
   U979 : NOR2_X1 port map( A1 => n425, A2 => n426, ZN => n298);
   U980 : NAND2_X1 port map( A1 => n603, A2 => n602, ZN => n393);
   U981 : INV_X1 port map( A => n407, ZN => n893);
   U982 : NAND2_X1 port map( A1 => n654, A2 => n655, ZN => n332);
   U983 : NAND2_X1 port map( A1 => n383, A2 => n384, ZN => n380);
   U984 : NAND2_X1 port map( A1 => n223, A2 => n224, ZN => n220);
   U985 : NAND2_X1 port map( A1 => n493, A2 => n494, ZN => n490);
   U986 : NAND2_X1 port map( A1 => n349, A2 => n348, ZN => n346);
   U987 : NAND2_X1 port map( A1 => n590, A2 => n580, ZN => n289);
   U988 : OAI211_X1 port map( C1 => n581, C2 => n582, A => n311, B => n310, ZN 
                           => n590);
   U989 : OR2_X1 port map( A1 => n589, A2 => n588, ZN => n583);
   U990 : NAND2_X1 port map( A1 => n587, A2 => n580, ZN => n288);
   U991 : OAI22_X1 port map( A1 => n581, A2 => n582, B1 => n310, B2 => n311, ZN
                           => n587);
   U992 : INV_X1 port map( A => n95, ZN => n950);
   U993 : INV_X1 port map( A => n166, ZN => n957);
   U994 : INV_X1 port map( A => n79, ZN => n948);
   U995 : INV_X1 port map( A => n87, ZN => n949);
   U996 : INV_X1 port map( A => n118, ZN => n951);
   U997 : INV_X1 port map( A => n126, ZN => n952);
   U998 : INV_X1 port map( A => n134, ZN => n953);
   U999 : INV_X1 port map( A => n142, ZN => n954);
   U1000 : INV_X1 port map( A => n150, ZN => n955);
   U1001 : INV_X1 port map( A => n158, ZN => n956);
   U1002 : INV_X1 port map( A => n176, ZN => n838);
   U1003 : NAND2_X1 port map( A1 => n588, A2 => n589, ZN => n584);
   U1004 : BUF_X1 port map( A => n47, Z => n800);
   U1005 : BUF_X1 port map( A => n47, Z => n801);
   U1006 : BUF_X1 port map( A => n47, Z => n802);
   U1007 : INV_X1 port map( A => n204, ZN => n943);
   U1008 : INV_X1 port map( A => n211, ZN => n941);
   U1009 : INV_X1 port map( A => n208, ZN => n942);
   U1010 : BUF_X1 port map( A => n185, Z => n797);
   U1011 : BUF_X1 port map( A => n185, Z => n798);
   U1012 : BUF_X1 port map( A => n185, Z => n799);
   U1013 : NAND4_X1 port map( A1 => n864, A2 => n863, A3 => n865, A4 => n665, 
                           ZN => n27);
   U1014 : NOR2_X1 port map( A1 => n663, A2 => n860, ZN => n665);
   U1015 : BUF_X1 port map( A => n778, Z => n795);
   U1016 : BUF_X1 port map( A => n778, Z => n791);
   U1017 : BUF_X1 port map( A => n778, Z => n792);
   U1018 : BUF_X1 port map( A => n778, Z => n790);
   U1019 : BUF_X1 port map( A => n778, Z => n793);
   U1020 : BUF_X1 port map( A => n778, Z => n794);
   U1021 : INV_X1 port map( A => n36, ZN => n841);
   U1022 : BUF_X1 port map( A => n778, Z => n796);
   U1023 : XNOR2_X1 port map( A => n783, B => RF_RD2_DATA(17), ZN => n459);
   U1024 : XNOR2_X1 port map( A => n785, B => RF_RD1_DATA(17), ZN => n458);
   U1025 : XNOR2_X1 port map( A => n785, B => RF_RD1_DATA(0), ZN => n426);
   U1026 : NAND4_X1 port map( A1 => n701, A2 => n699, A3 => n700, A4 => n947, 
                           ZN => n656);
   U1027 : OAI221_X1 port map( B1 => n900, B2 => n361, C1 => n362, C2 => n929, 
                           A => n364, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_24_port);
   U1028 : NAND2_X1 port map( A1 => n794, A2 => n929, ZN => n361);
   U1029 : AOI221_X1 port map( B1 => n791, B2 => n900, C1 => RF_RD1_DATA(24), 
                           C2 => n942, A => n941, ZN => n362);
   U1030 : AOI22_X1 port map( A1 => n365, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN291, B2 => n798, ZN => 
                           n364);
   U1031 : OAI221_X1 port map( B1 => n904, B2 => n411, C1 => n412, C2 => n931, 
                           A => n414, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_20_port);
   U1032 : NAND2_X1 port map( A1 => n794, A2 => n931, ZN => n411);
   U1033 : INV_X1 port map( A => RF_RD2_DATA(20), ZN => n931);
   U1034 : AOI221_X1 port map( B1 => n791, B2 => n904, C1 => RF_RD1_DATA(20), 
                           C2 => n942, A => n941, ZN => n412);
   U1035 : OAI221_X1 port map( B1 => n896, B2 => n314, C1 => n315, C2 => n927, 
                           A => n317, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_28_port);
   U1036 : NAND2_X1 port map( A1 => n793, A2 => n927, ZN => n314);
   U1037 : INV_X1 port map( A => RF_RD2_DATA(28), ZN => n927);
   U1038 : AOI221_X1 port map( B1 => n792, B2 => n896, C1 => RF_RD1_DATA(28), 
                           C2 => n942, A => n941, ZN => n315);
   U1039 : OAI221_X1 port map( B1 => n908, B2 => n471, C1 => n472, C2 => n933, 
                           A => n474, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_16_port);
   U1040 : NAND2_X1 port map( A1 => n794, A2 => n933, ZN => n471);
   U1041 : AOI221_X1 port map( B1 => n790, B2 => n908, C1 => RF_RD1_DATA(16), 
                           C2 => n942, A => n941, ZN => n472);
   U1042 : AOI22_X1 port map( A1 => n475, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN283, B2 => n797, ZN => 
                           n474);
   U1043 : NOR2_X1 port map( A1 => n947, A2 => n701, ZN => n564);
   U1044 : BUF_X1 port map( A => RF_RD2_DATA(3), Z => n816);
   U1045 : BUF_X1 port map( A => RF_RD2_DATA(2), Z => n818);
   U1046 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(13), ZN => n618);
   U1047 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(9), ZN => n627);
   U1048 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(9), ZN => n626);
   U1049 : XNOR2_X1 port map( A => n785, B => RF_RD1_DATA(1), ZN => n644);
   U1050 : XNOR2_X1 port map( A => n785, B => RF_RD1_DATA(5), ZN => n634);
   U1051 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(13), ZN => n617);
   U1052 : XNOR2_X1 port map( A => n783, B => RF_RD2_DATA(18), ZN => n652);
   U1053 : OAI211_X1 port map( C1 => n302, C2 => n926, A => n304, B => n305, ZN
                           => DATAPATH_IxThird_stxALU_out_i_29_port);
   U1054 : AOI221_X1 port map( B1 => n792, B2 => n895, C1 => RF_RD1_DATA(29), 
                           C2 => n942, A => n941, ZN => n302);
   U1055 : AOI22_X1 port map( A1 => n306, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN296, B2 => n798, ZN => 
                           n305);
   U1056 : NAND4_X1 port map( A1 => n700, A2 => n564, A3 => n565, A4 => n944, 
                           ZN => n552);
   U1057 : AOI21_X1 port map( B1 => n866, B2 => n573, A => n571, ZN => n566);
   U1058 : OAI211_X1 port map( C1 => n460, C2 => n932, A => n462, B => n463, ZN
                           => DATAPATH_IxThird_stxALU_out_i_17_port);
   U1059 : AOI221_X1 port map( B1 => n790, B2 => n907, C1 => RF_RD1_DATA(17), 
                           C2 => n942, A => n941, ZN => n460);
   U1060 : AOI22_X1 port map( A1 => n943, A2 => n464, B1 => 
                           DATAPATH_IxThird_stxALU1xN284, B2 => n797, ZN => 
                           n463);
   U1061 : OAI211_X1 port map( C1 => n320, C2 => n204, A => n321, B => n322, ZN
                           => DATAPATH_IxThird_stxALU_out_i_27_port);
   U1062 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(27), A3 => n897, ZN 
                           => n321);
   U1063 : AOI22_X1 port map( A1 => RF_RD2_DATA(27), A2 => n323, B1 => 
                           DATAPATH_IxThird_stxALU1xN294, B2 => n798, ZN => 
                           n322);
   U1064 : AOI22_X1 port map( A1 => n325, A2 => n326, B1 => n327, B2 => n869, 
                           ZN => n320);
   U1065 : OAI211_X1 port map( C1 => n336, C2 => n204, A => n337, B => n338, ZN
                           => DATAPATH_IxThird_stxALU_out_i_26_port);
   U1066 : OR3_X1 port map( A1 => n789, A2 => RF_RD2_DATA(26), A3 => n898, ZN 
                           => n337);
   U1067 : AOI22_X1 port map( A1 => RF_RD2_DATA(26), A2 => n339, B1 => 
                           DATAPATH_IxThird_stxALU1xN293, B2 => n798, ZN => 
                           n338);
   U1068 : AOI22_X1 port map( A1 => n341, A2 => n326, B1 => n342, B2 => n869, 
                           ZN => n336);
   U1069 : OAI211_X1 port map( C1 => n367, C2 => n204, A => n368, B => n369, ZN
                           => DATAPATH_IxThird_stxALU_out_i_23_port);
   U1070 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(23), A3 => n901, ZN 
                           => n368);
   U1071 : AOI22_X1 port map( A1 => RF_RD2_DATA(23), A2 => n370, B1 => 
                           DATAPATH_IxThird_stxALU1xN290, B2 => n798, ZN => 
                           n369);
   U1072 : AOI22_X1 port map( A1 => n372, A2 => n373, B1 => n870, B2 => n375, 
                           ZN => n367);
   U1073 : OAI211_X1 port map( C1 => n385, C2 => n204, A => n386, B => n387, ZN
                           => DATAPATH_IxThird_stxALU_out_i_22_port);
   U1074 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(22), A3 => n902, ZN 
                           => n386);
   U1075 : AOI22_X1 port map( A1 => RF_RD2_DATA(22), A2 => n388, B1 => 
                           DATAPATH_IxThird_stxALU1xN289, B2 => n798, ZN => 
                           n387);
   U1076 : AOI22_X1 port map( A1 => n390, A2 => n373, B1 => n391, B2 => n870, 
                           ZN => n385);
   U1077 : OAI211_X1 port map( C1 => n278, C2 => n204, A => n279, B => n280, ZN
                           => DATAPATH_IxThird_stxALU_out_i_30_port);
   U1078 : OR3_X1 port map( A1 => n789, A2 => RF_RD2_DATA(30), A3 => n894, ZN 
                           => n279);
   U1079 : AOI22_X1 port map( A1 => RF_RD2_DATA(30), A2 => n281, B1 => 
                           DATAPATH_IxThird_stxALU1xN297, B2 => n798, ZN => 
                           n280);
   U1080 : AOI22_X1 port map( A1 => n283, A2 => n866, B1 => n285, B2 => n286, 
                           ZN => n278);
   U1081 : OAI211_X1 port map( C1 => n428, C2 => n204, A => n429, B => n430, ZN
                           => DATAPATH_IxThird_stxALU_out_i_19_port);
   U1082 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(19), A3 => n905, ZN 
                           => n429);
   U1083 : AOI22_X1 port map( A1 => RF_RD2_DATA(19), A2 => n431, B1 => 
                           DATAPATH_IxThird_stxALU1xN286, B2 => n797, ZN => 
                           n430);
   U1084 : AOI22_X1 port map( A1 => n433, A2 => n876, B1 => n435, B2 => n436, 
                           ZN => n428);
   U1085 : OAI211_X1 port map( C1 => n444, C2 => n204, A => n445, B => n446, ZN
                           => DATAPATH_IxThird_stxALU_out_i_18_port);
   U1086 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(18), A3 => n906, ZN 
                           => n445);
   U1087 : AOI22_X1 port map( A1 => RF_RD2_DATA(18), A2 => n447, B1 => 
                           DATAPATH_IxThird_stxALU1xN285, B2 => n797, ZN => 
                           n446);
   U1088 : AOI22_X1 port map( A1 => n449, A2 => n876, B1 => n450, B2 => n436, 
                           ZN => n444);
   U1089 : OAI211_X1 port map( C1 => n350, C2 => n928, A => n352, B => n353, ZN
                           => DATAPATH_IxThird_stxALU_out_i_25_port);
   U1090 : AOI221_X1 port map( B1 => n791, B2 => n899, C1 => RF_RD1_DATA(25), 
                           C2 => n942, A => n941, ZN => n350);
   U1091 : AOI22_X1 port map( A1 => n943, A2 => n354, B1 => 
                           DATAPATH_IxThird_stxALU1xN292, B2 => n798, ZN => 
                           n353);
   U1092 : OAI211_X1 port map( C1 => n400, C2 => n930, A => n402, B => n403, ZN
                           => DATAPATH_IxThird_stxALU_out_i_21_port);
   U1093 : AOI221_X1 port map( B1 => n791, B2 => n903, C1 => RF_RD1_DATA(21), 
                           C2 => n942, A => n941, ZN => n400);
   U1094 : AOI22_X1 port map( A1 => n943, A2 => n404, B1 => 
                           DATAPATH_IxThird_stxALU1xN288, B2 => n798, ZN => 
                           n403);
   U1095 : INV_X1 port map( A => RF_RD1_DATA(6), ZN => n918);
   U1096 : INV_X1 port map( A => RF_RD1_DATA(2), ZN => n922);
   U1097 : INV_X1 port map( A => RF_RD1_DATA(10), ZN => n914);
   U1098 : INV_X1 port map( A => RF_RD2_DATA(8), ZN => n937);
   U1099 : INV_X1 port map( A => RF_RD2_DATA(4), ZN => n815);
   U1100 : INV_X1 port map( A => RF_RD1_DATA(4), ZN => n920);
   U1101 : INV_X1 port map( A => RF_RD1_DATA(8), ZN => n916);
   U1102 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(28), ZN => n311);
   U1103 : NOR3_X1 port map( A1 => n734, A2 => n733, A3 => n951, ZN => n109);
   U1104 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(28), ZN => n310);
   U1105 : INV_X1 port map( A => Rst, ZN => n840);
   U1106 : NOR3_X1 port map( A1 => n738, A2 => n737, A3 => n100, ZN => n95);
   U1107 : NOR3_X1 port map( A1 => n719, A2 => n718, A3 => n720, ZN => n166);
   U1108 : NOR3_X1 port map( A1 => n742, A2 => n741, A3 => n949, ZN => n79);
   U1109 : NOR3_X1 port map( A1 => n740, A2 => n739, A3 => n950, ZN => n87);
   U1110 : NOR3_X1 port map( A1 => n732, A2 => n731, A3 => n952, ZN => n118);
   U1111 : NOR3_X1 port map( A1 => n730, A2 => n729, A3 => n953, ZN => n126);
   U1112 : NOR3_X1 port map( A1 => n728, A2 => n727, A3 => n954, ZN => n134);
   U1113 : NOR3_X1 port map( A1 => n726, A2 => n725, A3 => n955, ZN => n142);
   U1114 : NOR3_X1 port map( A1 => n724, A2 => n723, A3 => n956, ZN => n150);
   U1115 : NOR3_X1 port map( A1 => n722, A2 => n721, A3 => n957, ZN => n158);
   U1116 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(29), ZN => n581);
   U1117 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(25), ZN => n349);
   U1118 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(25), ZN => n348);
   U1119 : NOR3_X1 port map( A1 => n744, A2 => n743, A3 => n948, ZN => n72);
   U1120 : AOI21_X1 port map( B1 => n804, B2 => n718, A => n83, ZN => n176);
   U1121 : OAI221_X1 port map( B1 => n912, B2 => n518, C1 => n519, C2 => n935, 
                           A => n521, ZN => 
                           DATAPATH_IxThird_stxALU_out_i_12_port);
   U1122 : NAND2_X1 port map( A1 => n794, A2 => n935, ZN => n518);
   U1123 : AOI221_X1 port map( B1 => n790, B2 => n912, C1 => RF_RD1_DATA(12), 
                           C2 => n942, A => n941, ZN => n519);
   U1124 : AOI22_X1 port map( A1 => n522, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN279, B2 => n797, ZN => 
                           n521);
   U1125 : AND2_X1 port map( A1 => n72, A2 => IRAM_ADD_29_port, ZN => n65);
   U1126 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(21), ZN => n602);
   U1127 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(21), ZN => n603);
   U1128 : OAI22_X1 port map( A1 => n718, A2 => n839, B1 => n810, B2 => 
                           IRAM_ADD_2_port, ZN => n777);
   U1129 : OAI22_X1 port map( A1 => n703, A2 => n839, B1 => n811, B2 => n859, 
                           ZN => n682);
   U1130 : INV_X1 port map( A => IRAM_DOUT(7), ZN => n859);
   U1131 : OAI22_X1 port map( A1 => n704, A2 => n839, B1 => n811, B2 => n858, 
                           ZN => n683);
   U1132 : INV_X1 port map( A => IRAM_DOUT(8), ZN => n858);
   U1133 : OAI22_X1 port map( A1 => n705, A2 => n839, B1 => n810, B2 => n857, 
                           ZN => n684);
   U1134 : INV_X1 port map( A => IRAM_DOUT(9), ZN => n857);
   U1135 : OAI22_X1 port map( A1 => n706, A2 => n839, B1 => n811, B2 => n856, 
                           ZN => n685);
   U1136 : INV_X1 port map( A => IRAM_DOUT(10), ZN => n856);
   U1137 : OAI22_X1 port map( A1 => n707, A2 => n839, B1 => n808, B2 => n855, 
                           ZN => n686);
   U1138 : INV_X1 port map( A => IRAM_DOUT(11), ZN => n855);
   U1139 : OAI22_X1 port map( A1 => n708, A2 => n839, B1 => n810, B2 => n851, 
                           ZN => n687);
   U1140 : INV_X1 port map( A => IRAM_DOUT(15), ZN => n851);
   U1141 : OAI22_X1 port map( A1 => n709, A2 => n839, B1 => n810, B2 => n850, 
                           ZN => n688);
   U1142 : INV_X1 port map( A => IRAM_DOUT(16), ZN => n850);
   U1143 : OAI22_X1 port map( A1 => n710, A2 => n839, B1 => n809, B2 => n849, 
                           ZN => n689);
   U1144 : INV_X1 port map( A => IRAM_DOUT(17), ZN => n849);
   U1145 : OAI22_X1 port map( A1 => n711, A2 => n839, B1 => n809, B2 => n848, 
                           ZN => n690);
   U1146 : INV_X1 port map( A => IRAM_DOUT(18), ZN => n848);
   U1147 : OAI22_X1 port map( A1 => n712, A2 => n839, B1 => n809, B2 => n847, 
                           ZN => n691);
   U1148 : INV_X1 port map( A => IRAM_DOUT(19), ZN => n847);
   U1149 : OAI22_X1 port map( A1 => n713, A2 => n839, B1 => n809, B2 => n846, 
                           ZN => n692);
   U1150 : INV_X1 port map( A => IRAM_DOUT(20), ZN => n846);
   U1151 : OAI22_X1 port map( A1 => n714, A2 => n839, B1 => n808, B2 => n845, 
                           ZN => n693);
   U1152 : INV_X1 port map( A => IRAM_DOUT(21), ZN => n845);
   U1153 : OAI22_X1 port map( A1 => n715, A2 => n839, B1 => n808, B2 => n844, 
                           ZN => n694);
   U1154 : INV_X1 port map( A => IRAM_DOUT(22), ZN => n844);
   U1155 : OAI22_X1 port map( A1 => n716, A2 => n839, B1 => n808, B2 => n843, 
                           ZN => n695);
   U1156 : INV_X1 port map( A => IRAM_DOUT(23), ZN => n843);
   U1157 : OAI22_X1 port map( A1 => n717, A2 => n839, B1 => n807, B2 => n842, 
                           ZN => n696);
   U1158 : INV_X1 port map( A => IRAM_DOUT(24), ZN => n842);
   U1159 : OAI211_X1 port map( C1 => n247, C2 => n815, A => n249, B => n250, ZN
                           => DATAPATH_IxThird_stxALU_out_i_4_port);
   U1160 : AOI221_X1 port map( B1 => n792, B2 => n920, C1 => RF_RD1_DATA(4), C2
                           => n942, A => n941, ZN => n247);
   U1161 : AOI22_X1 port map( A1 => n251, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN271, B2 => n799, ZN => 
                           n250);
   U1162 : OAI211_X1 port map( C1 => n196, C2 => n937, A => n198, B => n199, ZN
                           => DATAPATH_IxThird_stxALU_out_i_8_port);
   U1163 : AOI221_X1 port map( B1 => n793, B2 => n916, C1 => RF_RD1_DATA(8), C2
                           => n942, A => n941, ZN => n196);
   U1164 : AOI22_X1 port map( A1 => n200, A2 => n943, B1 => 
                           DATAPATH_IxThird_stxALU1xN275, B2 => n799, ZN => 
                           n199);
   U1165 : OAI211_X1 port map( C1 => n179, C2 => n936, A => n181, B => n182, ZN
                           => DATAPATH_IxThird_stxALU_out_i_9_port);
   U1166 : AOI221_X1 port map( B1 => n793, B2 => n915, C1 => n942, C2 => 
                           RF_RD1_DATA(9), A => n941, ZN => n179);
   U1167 : AOI22_X1 port map( A1 => n943, A2 => n184, B1 => 
                           DATAPATH_IxThird_stxALU1xN276, B2 => n799, ZN => 
                           n182);
   U1168 : OAI211_X1 port map( C1 => n477, C2 => n204, A => n478, B => n479, ZN
                           => DATAPATH_IxThird_stxALU_out_i_15_port);
   U1169 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(15), A3 => n909, ZN 
                           => n478);
   U1170 : AOI22_X1 port map( A1 => RF_RD2_DATA(15), A2 => n480, B1 => 
                           DATAPATH_IxThird_stxALU1xN282, B2 => n797, ZN => 
                           n479);
   U1171 : AOI22_X1 port map( A1 => n482, A2 => n483, B1 => n878, B2 => n485, 
                           ZN => n477);
   U1172 : OAI211_X1 port map( C1 => n495, C2 => n204, A => n496, B => n497, ZN
                           => DATAPATH_IxThird_stxALU_out_i_14_port);
   U1173 : OR3_X1 port map( A1 => n789, A2 => RF_RD2_DATA(14), A3 => n910, ZN 
                           => n496);
   U1174 : AOI22_X1 port map( A1 => RF_RD2_DATA(14), A2 => n498, B1 => 
                           DATAPATH_IxThird_stxALU1xN281, B2 => n797, ZN => 
                           n497);
   U1175 : AOI22_X1 port map( A1 => n500, A2 => n483, B1 => n501, B2 => n878, 
                           ZN => n495);
   U1176 : OAI211_X1 port map( C1 => n507, C2 => n934, A => n509, B => n510, ZN
                           => DATAPATH_IxThird_stxALU_out_i_13_port);
   U1177 : AOI221_X1 port map( B1 => n790, B2 => n911, C1 => RF_RD1_DATA(13), 
                           C2 => n942, A => n941, ZN => n507);
   U1178 : AOI22_X1 port map( A1 => n943, A2 => n511, B1 => 
                           DATAPATH_IxThird_stxALU1xN280, B2 => n797, ZN => 
                           n510);
   U1179 : OAI211_X1 port map( C1 => n524, C2 => n204, A => n525, B => n526, ZN
                           => DATAPATH_IxThird_stxALU_out_i_11_port);
   U1180 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(11), A3 => n913, ZN 
                           => n525);
   U1181 : AOI22_X1 port map( A1 => RF_RD2_DATA(11), A2 => n527, B1 => 
                           DATAPATH_IxThird_stxALU1xN278, B2 => n797, ZN => 
                           n526);
   U1182 : AOI22_X1 port map( A1 => n529, A2 => n882, B1 => n531, B2 => n191, 
                           ZN => n524);
   U1183 : OAI211_X1 port map( C1 => n225, C2 => n204, A => n226, B => n227, ZN
                           => DATAPATH_IxThird_stxALU_out_i_6_port);
   U1184 : OR3_X1 port map( A1 => n789, A2 => RF_RD2_DATA(6), A3 => n918, ZN =>
                           n226);
   U1185 : AOI22_X1 port map( A1 => RF_RD2_DATA(6), A2 => n228, B1 => 
                           DATAPATH_IxThird_stxALU1xN273, B2 => n799, ZN => 
                           n227);
   U1186 : AOI22_X1 port map( A1 => n230, A2 => n884, B1 => n231, B2 => n215, 
                           ZN => n225);
   U1187 : OAI211_X1 port map( C1 => n539, C2 => n204, A => n540, B => n541, ZN
                           => DATAPATH_IxThird_stxALU_out_i_10_port);
   U1188 : OR3_X1 port map( A1 => n789, A2 => RF_RD2_DATA(10), A3 => n914, ZN 
                           => n540);
   U1189 : AOI22_X1 port map( A1 => RF_RD2_DATA(10), A2 => n542, B1 => 
                           DATAPATH_IxThird_stxALU1xN277, B2 => n797, ZN => 
                           n541);
   U1190 : AOI22_X1 port map( A1 => n544, A2 => n882, B1 => n545, B2 => n191, 
                           ZN => n539);
   U1191 : OAI211_X1 port map( C1 => n203, C2 => n204, A => n205, B => n206, ZN
                           => DATAPATH_IxThird_stxALU_out_i_7_port);
   U1192 : OR3_X1 port map( A1 => n788, A2 => RF_RD2_DATA(7), A3 => n917, ZN =>
                           n205);
   U1193 : AOI22_X1 port map( A1 => RF_RD2_DATA(7), A2 => n207, B1 => 
                           DATAPATH_IxThird_stxALU1xN274, B2 => n799, ZN => 
                           n206);
   U1194 : AOI22_X1 port map( A1 => n884, A2 => n213, B1 => n214, B2 => n215, 
                           ZN => n203);
   U1195 : XNOR2_X1 port map( A => n782, B => RF_RD2_DATA(30), ZN => n589);
   U1196 : XNOR2_X1 port map( A => n786, B => RF_RD1_DATA(30), ZN => n588);
   U1197 : OAI21_X1 port map( B1 => n745, B2 => n73, A => n74, ZN => n750);
   U1198 : AOI21_X1 port map( B1 => n744, B2 => n803, A => n76, ZN => n73);
   U1199 : OAI21_X1 port map( B1 => n736, B2 => n110, A => n111, ZN => n759);
   U1200 : NAND4_X1 port map( A1 => n736, A2 => n109, A3 => n803, A4 => 
                           IRAM_ADD_19_port, ZN => n111);
   U1201 : AOI21_X1 port map( B1 => n735, B2 => n804, A => n112, ZN => n110);
   U1202 : NAND2_X1 port map( A1 => Rst, A2 => n839, ZN => n47);
   U1203 : BUF_X1 port map( A => RF_RD2_DATA(0), Z => n823);
   U1204 : OAI22_X1 port map( A1 => n738, A2 => n101, B1 => n83, B2 => n102, ZN
                           => n757);
   U1205 : NOR3_X1 port map( A1 => n100, A2 => n737, A3 => n83, ZN => n101);
   U1206 : AOI21_X1 port map( B1 => n103, B2 => n738, A => n840, ZN => n102);
   U1207 : NOR2_X1 port map( A1 => n737, A2 => n100, ZN => n103);
   U1208 : OAI21_X1 port map( B1 => n734, B2 => n831, A => n117, ZN => n761);
   U1209 : NAND4_X1 port map( A1 => n734, A2 => n118, A3 => n803, A4 => 
                           IRAM_ADD_17_port, ZN => n117);
   U1210 : INV_X1 port map( A => n120, ZN => n831);
   U1211 : OAI21_X1 port map( B1 => IRAM_ADD_17_port, B2 => n806, A => n121, ZN
                           => n120);
   U1212 : OAI21_X1 port map( B1 => n732, B2 => n832, A => n125, ZN => n763);
   U1213 : NAND4_X1 port map( A1 => n732, A2 => n126, A3 => n803, A4 => 
                           IRAM_ADD_15_port, ZN => n125);
   U1214 : INV_X1 port map( A => n128, ZN => n832);
   U1215 : OAI21_X1 port map( B1 => IRAM_ADD_15_port, B2 => n806, A => n129, ZN
                           => n128);
   U1216 : OAI21_X1 port map( B1 => n730, B2 => n833, A => n133, ZN => n765);
   U1217 : NAND4_X1 port map( A1 => n730, A2 => n134, A3 => n803, A4 => 
                           IRAM_ADD_13_port, ZN => n133);
   U1218 : INV_X1 port map( A => n136, ZN => n833);
   U1219 : OAI21_X1 port map( B1 => IRAM_ADD_13_port, B2 => n806, A => n137, ZN
                           => n136);
   U1220 : OAI21_X1 port map( B1 => n728, B2 => n834, A => n141, ZN => n767);
   U1221 : NAND4_X1 port map( A1 => n728, A2 => n142, A3 => n803, A4 => 
                           IRAM_ADD_11_port, ZN => n141);
   U1222 : INV_X1 port map( A => n144, ZN => n834);
   U1223 : OAI21_X1 port map( B1 => IRAM_ADD_11_port, B2 => n805, A => n145, ZN
                           => n144);
   U1224 : OAI21_X1 port map( B1 => n726, B2 => n835, A => n149, ZN => n769);
   U1225 : NAND4_X1 port map( A1 => n726, A2 => n150, A3 => n803, A4 => 
                           IRAM_ADD_9_port, ZN => n149);
   U1226 : INV_X1 port map( A => n152, ZN => n835);
   U1227 : OAI21_X1 port map( B1 => IRAM_ADD_9_port, B2 => n805, A => n153, ZN 
                           => n152);
   U1228 : OAI21_X1 port map( B1 => n724, B2 => n836, A => n157, ZN => n771);
   U1229 : NAND4_X1 port map( A1 => n724, A2 => n158, A3 => n803, A4 => 
                           IRAM_ADD_7_port, ZN => n157);
   U1230 : INV_X1 port map( A => n160, ZN => n836);
   U1231 : OAI21_X1 port map( B1 => IRAM_ADD_7_port, B2 => n805, A => n161, ZN 
                           => n160);
   U1232 : OAI21_X1 port map( B1 => n722, B2 => n837, A => n165, ZN => n773);
   U1233 : NAND4_X1 port map( A1 => n722, A2 => n166, A3 => n803, A4 => 
                           IRAM_ADD_5_port, ZN => n165);
   U1234 : INV_X1 port map( A => n168, ZN => n837);
   U1235 : OAI21_X1 port map( B1 => IRAM_ADD_5_port, B2 => n805, A => n169, ZN 
                           => n168);
   U1236 : OAI21_X1 port map( B1 => n742, B2 => n829, A => n86, ZN => n753);
   U1237 : NAND4_X1 port map( A1 => n742, A2 => n87, A3 => n804, A4 => 
                           IRAM_ADD_25_port, ZN => n86);
   U1238 : INV_X1 port map( A => n89, ZN => n829);
   U1239 : OAI21_X1 port map( B1 => IRAM_ADD_25_port, B2 => n807, A => n90, ZN 
                           => n89);
   U1240 : OAI21_X1 port map( B1 => n740, B2 => n830, A => n94, ZN => n755);
   U1241 : NAND4_X1 port map( A1 => n740, A2 => n95, A3 => n803, A4 => 
                           IRAM_ADD_23_port, ZN => n94);
   U1242 : INV_X1 port map( A => n97, ZN => n830);
   U1243 : OAI21_X1 port map( B1 => IRAM_ADD_23_port, B2 => n807, A => n98, ZN 
                           => n97);
   U1244 : OAI211_X1 port map( C1 => n237, C2 => n814, A => n239, B => n240, ZN
                           => DATAPATH_IxThird_stxALU_out_i_5_port);
   U1245 : AOI221_X1 port map( B1 => n793, B2 => n919, C1 => RF_RD1_DATA(5), C2
                           => n942, A => n941, ZN => n237);
   U1246 : AOI22_X1 port map( A1 => n943, A2 => n241, B1 => 
                           DATAPATH_IxThird_stxALU1xN272, B2 => n799, ZN => 
                           n240);
   U1247 : INV_X1 port map( A => RF_RD1_DATA(22), ZN => n902);
   U1248 : INV_X1 port map( A => RF_RD1_DATA(14), ZN => n910);
   U1249 : OAI21_X1 port map( B1 => n719, B2 => n176, A => n177, ZN => n776);
   U1250 : OAI21_X1 port map( B1 => n743, B2 => n81, A => n82, ZN => n752);
   U1251 : OAI21_X1 port map( B1 => n741, B2 => n90, A => n91, ZN => n754);
   U1252 : OAI21_X1 port map( B1 => n739, B2 => n98, A => n99, ZN => n756);
   U1253 : OAI21_X1 port map( B1 => n733, B2 => n121, A => n122, ZN => n762);
   U1254 : OAI21_X1 port map( B1 => n731, B2 => n129, A => n130, ZN => n764);
   U1255 : OAI21_X1 port map( B1 => n729, B2 => n137, A => n138, ZN => n766);
   U1256 : OAI21_X1 port map( B1 => n727, B2 => n145, A => n146, ZN => n768);
   U1257 : OAI21_X1 port map( B1 => n725, B2 => n153, A => n154, ZN => n770);
   U1258 : OAI21_X1 port map( B1 => n723, B2 => n161, A => n162, ZN => n772);
   U1259 : OAI21_X1 port map( B1 => n721, B2 => n169, A => n170, ZN => n774);
   U1260 : OAI21_X1 port map( B1 => n746, B2 => n826, A => n70, ZN => n749);
   U1261 : INV_X1 port map( A => n68, ZN => n826);
   U1262 : OAI21_X1 port map( B1 => n735, B2 => n827, A => n114, ZN => n760);
   U1263 : INV_X1 port map( A => n112, ZN => n827);
   U1264 : OAI21_X1 port map( B1 => n720, B2 => n171, A => n172, ZN => n775);
   U1265 : NAND4_X1 port map( A1 => n720, A2 => n804, A3 => IRAM_ADD_3_port, A4
                           => IRAM_ADD_2_port, ZN => n172);
   U1266 : AOI21_X1 port map( B1 => n719, B2 => n803, A => n838, ZN => n171);
   U1267 : INV_X1 port map( A => RF_RD2_DATA(31), ZN => n925);
   U1268 : OAI21_X1 port map( B1 => n747, B2 => n63, A => n64, ZN => n748);
   U1269 : NAND4_X1 port map( A1 => n747, A2 => n65, A3 => n803, A4 => 
                           IRAM_ADD_30_port, ZN => n64);
   U1270 : AOI21_X1 port map( B1 => n746, B2 => n804, A => n68, ZN => n63);
   U1271 : INV_X1 port map( A => RF_RD2_DATA(24), ZN => n929);
   U1272 : INV_X1 port map( A => RF_RD2_DATA(16), ZN => n933);
   U1273 : INV_X1 port map( A => RF_RD2_DATA(12), ZN => n935);
   U1274 : INV_X1 port map( A => RF_RD1_DATA(24), ZN => n900);
   U1275 : INV_X1 port map( A => RF_RD1_DATA(16), ZN => n908);
   U1276 : INV_X1 port map( A => RF_RD1_DATA(20), ZN => n904);
   U1277 : INV_X1 port map( A => RF_RD1_DATA(12), ZN => n912);
   U1278 : INV_X1 port map( A => RF_RD1_DATA(18), ZN => n906);
   U1279 : INV_X1 port map( A => RF_RD2_DATA(29), ZN => n926);
   U1280 : OAI22_X1 port map( A1 => n737, A2 => n104, B1 => IRAM_ADD_21_port, 
                           B2 => n106, ZN => n758);
   U1281 : AOI21_X1 port map( B1 => n804, B2 => n100, A => n83, ZN => n104);
   U1282 : OR2_X1 port map( A1 => n100, A2 => n812, ZN => n106);
   U1283 : OAI21_X1 port map( B1 => n744, B2 => n828, A => n78, ZN => n751);
   U1284 : NAND4_X1 port map( A1 => n744, A2 => n79, A3 => n804, A4 => 
                           IRAM_ADD_27_port, ZN => n78);
   U1285 : INV_X1 port map( A => n76, ZN => n828);
   U1286 : NAND4_X1 port map( A1 => n701, A2 => n702, A3 => n945, A4 => n944, 
                           ZN => n211);
   U1287 : NOR4_X1 port map( A1 => n854, A2 => n41, A3 => IRAM_DOUT(2), A4 => 
                           IRAM_DOUT(5), ZN => n36);
   U1288 : NAND3_X1 port map( A1 => n701, A2 => n702, A3 => n556, ZN => n208);
   U1289 : NOR3_X1 port map( A1 => n700, A2 => n699, A3 => n946, ZN => n185);
   U1290 : NOR2_X1 port map( A1 => n944, A2 => n700, ZN => n556);
   U1291 : OAI221_X1 port map( B1 => n208, B2 => n897, C1 => RF_RD1_DATA(27), 
                           C2 => n789, A => n211, ZN => n323);
   U1292 : OAI221_X1 port map( B1 => n208, B2 => n898, C1 => RF_RD1_DATA(26), 
                           C2 => n789, A => n211, ZN => n339);
   U1293 : OAI221_X1 port map( B1 => n208, B2 => n901, C1 => RF_RD1_DATA(23), 
                           C2 => n789, A => n211, ZN => n370);
   U1294 : OAI221_X1 port map( B1 => n208, B2 => n902, C1 => RF_RD1_DATA(22), 
                           C2 => n789, A => n211, ZN => n388);
   U1295 : OAI221_X1 port map( B1 => n208, B2 => n905, C1 => RF_RD1_DATA(19), 
                           C2 => n789, A => n211, ZN => n431);
   U1296 : OAI221_X1 port map( B1 => n208, B2 => n906, C1 => RF_RD1_DATA(18), 
                           C2 => n789, A => n211, ZN => n447);
   U1297 : OAI221_X1 port map( B1 => n208, B2 => n913, C1 => RF_RD1_DATA(11), 
                           C2 => n788, A => n211, ZN => n527);
   U1298 : OAI221_X1 port map( B1 => n208, B2 => n917, C1 => RF_RD1_DATA(7), C2
                           => n788, A => n211, ZN => n207);
   U1299 : OAI221_X1 port map( B1 => n208, B2 => n918, C1 => RF_RD1_DATA(6), C2
                           => n788, A => n211, ZN => n228);
   U1300 : OAI221_X1 port map( B1 => n208, B2 => n894, C1 => RF_RD1_DATA(30), 
                           C2 => n789, A => n211, ZN => n281);
   U1301 : OAI221_X1 port map( B1 => n208, B2 => n921, C1 => RF_RD1_DATA(3), C2
                           => n789, A => n211, ZN => n257);
   U1302 : OAI221_X1 port map( B1 => n208, B2 => n922, C1 => RF_RD1_DATA(2), C2
                           => n789, A => n211, ZN => n293);
   U1303 : OAI221_X1 port map( B1 => n208, B2 => n923, C1 => RF_RD1_DATA(1), C2
                           => n789, A => n211, ZN => n420);
   U1304 : OAI221_X1 port map( B1 => n208, B2 => n909, C1 => RF_RD1_DATA(15), 
                           C2 => n788, A => n211, ZN => n480);
   U1305 : OAI221_X1 port map( B1 => n208, B2 => n910, C1 => RF_RD1_DATA(14), 
                           C2 => n788, A => n211, ZN => n498);
   U1306 : OAI221_X1 port map( B1 => n208, B2 => n914, C1 => RF_RD1_DATA(10), 
                           C2 => n788, A => n211, ZN => n542);
   U1307 : OAI221_X1 port map( B1 => n208, B2 => n924, C1 => RF_RD1_DATA(0), C2
                           => n788, A => n211, ZN => n561);
   U1308 : AND3_X1 port map( A1 => n700, A2 => n564, A3 => n699, ZN => n778);
   U1309 : NOR2_X1 port map( A1 => n861, A2 => n41, ZN => n28);
   U1310 : INV_X1 port map( A => IRAM_DOUT(5), ZN => n861);
   U1311 : OAI22_X1 port map( A1 => n27, A2 => n840, B1 => Rst, B2 => n670, ZN 
                           => n26);
   U1312 : BUF_X1 port map( A => RF_RD2_DATA(3), Z => n817);
   U1313 : BUF_X1 port map( A => RF_RD2_DATA(2), Z => n819);
   U1314 : OAI22_X1 port map( A1 => n670, A2 => n840, B1 => n701, B2 => Rst, ZN
                           => n675);
   U1315 : OAI22_X1 port map( A1 => n671, A2 => n840, B1 => n700, B2 => Rst, ZN
                           => n676);
   U1316 : OAI22_X1 port map( A1 => n669, A2 => n840, B1 => n702, B2 => Rst, ZN
                           => n674);
   U1317 : OAI22_X1 port map( A1 => n672, A2 => n840, B1 => n699, B2 => Rst, ZN
                           => n677);
   U1318 : OAI22_X1 port map( A1 => n698, A2 => n939, B1 => n938, B2 => n27, ZN
                           => CU_IxN52);
   U1319 : INV_X1 port map( A => n659, ZN => n938);
   U1320 : OAI22_X1 port map( A1 => n669, A2 => Rst, B1 => n21, B2 => n841, ZN 
                           => n678);
   U1321 : INV_X1 port map( A => IRAM_DOUT(13), ZN => n853);
   U1322 : NAND4_X1 port map( A1 => n864, A2 => n860, A3 => Rst, A4 => n45, ZN 
                           => n41);
   U1323 : AND3_X1 port map( A1 => IRAM_DOUT(4), A2 => IRAM_DOUT(0), A3 => 
                           IRAM_DOUT(1), ZN => n45);
   U1324 : BUF_X1 port map( A => RF_RD2_DATA(1), Z => n821);
   U1325 : NAND2_X1 port map( A1 => IRAM_DOUT(13), A2 => n852, ZN => n21);
   U1326 : OAI211_X1 port map( C1 => n841, C2 => n852, A => n33, B => n825, ZN 
                           => n680);
   U1327 : INV_X1 port map( A => n35, ZN => n825);
   U1328 : OAI22_X1 port map( A1 => n27, A2 => n840, B1 => Rst, B2 => n671, ZN 
                           => n35);
   U1329 : INV_X1 port map( A => IRAM_DOUT(2), ZN => n865);
   U1330 : OAI21_X1 port map( B1 => n698, B2 => n939, A => n658, ZN => CU_IxN53
                           );
   U1331 : NAND4_X1 port map( A1 => n659, A2 => n863, A3 => n862, A4 => n662, 
                           ZN => n658);
   U1332 : INV_X1 port map( A => n663, ZN => n862);
   U1333 : NOR3_X1 port map( A1 => n864, A2 => n860, A3 => n865, ZN => n662);
   U1334 : INV_X1 port map( A => IRAM_DOUT(6), ZN => n860);
   U1335 : NAND2_X1 port map( A1 => n698, A2 => n939, ZN => n659);
   U1336 : INV_X1 port map( A => IRAM_DOUT(14), ZN => n852);
   U1337 : INV_X1 port map( A => IRAM_DOUT(3), ZN => n864);
   U1338 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n854, A4 => n865, ZN 
                           => n23);
   U1339 : INV_X1 port map( A => n26, ZN => n824);
   U1340 : OAI21_X1 port map( B1 => IRAM_DOUT(13), B2 => n852, A => n21, ZN => 
                           n29);
   U1341 : AOI22_X1 port map( A1 => n38, A2 => n28, B1 => n840, B2 => n940, ZN 
                           => n37);
   U1342 : NOR2_X1 port map( A1 => IRAM_DOUT(12), A2 => n21, ZN => n38);
   U1343 : NAND2_X1 port map( A1 => IRAM_DOUT(2), A2 => n28, ZN => n33);
   U1344 : NOR2_X1 port map( A1 => n667, A2 => n840, ZN => n697);
   U1345 : NOR2_X1 port map( A1 => n668, A2 => n840, ZN => n673);
   U1346 : INV_X1 port map( A => IRAM_DOUT(12), ZN => n854);
   U1347 : INV_X1 port map( A => RF_RD1_DATA(28), ZN => n896);
   U1348 : INV_X1 port map( A => IRAM_DOUT(4), ZN => n863);
   U1349 : INV_X1 port map( A => RF_RD1_DATA(27), ZN => n897);
   U1350 : INV_X1 port map( A => RF_RD1_DATA(26), ZN => n898);
   U1351 : INV_X1 port map( A => RF_RD1_DATA(23), ZN => n901);
   U1352 : INV_X1 port map( A => RF_RD1_DATA(19), ZN => n905);
   U1353 : INV_X1 port map( A => RF_RD1_DATA(11), ZN => n913);
   U1354 : INV_X1 port map( A => RF_RD1_DATA(7), ZN => n917);
   U1355 : INV_X1 port map( A => RF_RD1_DATA(30), ZN => n894);
   U1356 : INV_X1 port map( A => RF_RD1_DATA(3), ZN => n921);
   U1357 : INV_X1 port map( A => RF_RD1_DATA(1), ZN => n923);
   U1358 : INV_X1 port map( A => RF_RD1_DATA(15), ZN => n909);
   U1359 : INV_X1 port map( A => RF_RD1_DATA(0), ZN => n924);
   U1360 : INV_X1 port map( A => RF_RD2_DATA(25), ZN => n928);
   U1361 : INV_X1 port map( A => RF_RD2_DATA(21), ZN => n930);
   U1362 : INV_X1 port map( A => RF_RD2_DATA(13), ZN => n934);
   U1363 : INV_X1 port map( A => RF_RD2_DATA(9), ZN => n936);
   U1364 : INV_X1 port map( A => RF_RD2_DATA(17), ZN => n932);
   U1365 : INV_X1 port map( A => RF_RD1_DATA(25), ZN => n899);
   U1366 : INV_X1 port map( A => RF_RD1_DATA(21), ZN => n903);
   U1367 : INV_X1 port map( A => RF_RD1_DATA(13), ZN => n911);
   U1368 : INV_X1 port map( A => RF_RD1_DATA(5), ZN => n919);
   U1369 : INV_X1 port map( A => RF_RD1_DATA(29), ZN => n895);
   U1370 : INV_X1 port map( A => RF_RD1_DATA(9), ZN => n915);
   U1371 : INV_X1 port map( A => RF_RD1_DATA(17), ZN => n907);
   U1372 : INV_X1 port map( A => RF_RD1_DATA(31), ZN => n813);
   U1373 : INV_X1 port map( A => RF_RD2_DATA(5), ZN => n814);
   U1374 : MUX2_X1 port map( A => RF_RD1_DATA(0), B => RF_RD1_DATA(1), S => 
                           n822, Z => n958);
   U1375 : MUX2_X1 port map( A => RF_RD1_DATA(2), B => RF_RD1_DATA(3), S => 
                           n822, Z => n1054);
   U1376 : MUX2_X1 port map( A => n958, B => n1054, S => n820, Z => n959);
   U1377 : MUX2_X1 port map( A => RF_RD1_DATA(4), B => RF_RD1_DATA(5), S => 
                           n822, Z => n1053);
   U1378 : MUX2_X1 port map( A => RF_RD1_DATA(6), B => RF_RD1_DATA(7), S => 
                           n822, Z => n1056);
   U1379 : MUX2_X1 port map( A => n1053, B => n1056, S => n820, Z => n1076);
   U1380 : MUX2_X1 port map( A => n959, B => n1076, S => n818, Z => n960);
   U1381 : MUX2_X1 port map( A => RF_RD1_DATA(8), B => RF_RD1_DATA(9), S => 
                           n822, Z => n1055);
   U1382 : MUX2_X1 port map( A => RF_RD1_DATA(10), B => RF_RD1_DATA(11), S => 
                           n822, Z => n964);
   U1383 : MUX2_X1 port map( A => n1055, B => n964, S => n820, Z => n1075);
   U1384 : MUX2_X1 port map( A => RF_RD1_DATA(12), B => RF_RD1_DATA(13), S => 
                           n822, Z => n963);
   U1385 : MUX2_X1 port map( A => RF_RD1_DATA(14), B => RF_RD1_DATA(15), S => 
                           n822, Z => n966);
   U1386 : MUX2_X1 port map( A => n963, B => n966, S => n820, Z => n979);
   U1387 : MUX2_X1 port map( A => n1075, B => n979, S => n818, Z => n1104);
   U1388 : MUX2_X1 port map( A => n960, B => n1104, S => n816, Z => n961);
   U1389 : MUX2_X1 port map( A => RF_RD1_DATA(16), B => RF_RD1_DATA(17), S => 
                           n822, Z => n965);
   U1390 : MUX2_X1 port map( A => RF_RD1_DATA(18), B => RF_RD1_DATA(19), S => 
                           n822, Z => n968);
   U1391 : MUX2_X1 port map( A => n965, B => n968, S => n820, Z => n978);
   U1392 : MUX2_X1 port map( A => RF_RD1_DATA(20), B => RF_RD1_DATA(21), S => 
                           n822, Z => n967);
   U1393 : MUX2_X1 port map( A => RF_RD1_DATA(22), B => RF_RD1_DATA(23), S => 
                           n822, Z => n970);
   U1394 : MUX2_X1 port map( A => n967, B => n970, S => n820, Z => n981);
   U1395 : MUX2_X1 port map( A => n978, B => n981, S => n818, Z => n1103);
   U1396 : MUX2_X1 port map( A => RF_RD1_DATA(24), B => RF_RD1_DATA(25), S => 
                           n822, Z => n969);
   U1397 : MUX2_X1 port map( A => RF_RD1_DATA(26), B => RF_RD1_DATA(27), S => 
                           n822, Z => n972);
   U1398 : MUX2_X1 port map( A => n969, B => n972, S => n820, Z => n980);
   U1399 : MUX2_X1 port map( A => RF_RD1_DATA(28), B => RF_RD1_DATA(29), S => 
                           n822, Z => n971);
   U1400 : MUX2_X1 port map( A => RF_RD1_DATA(30), B => n781, S => n822, Z => 
                           n973);
   U1401 : MUX2_X1 port map( A => n971, B => n973, S => n820, Z => n982);
   U1402 : MUX2_X1 port map( A => n980, B => n982, S => n818, Z => n1041);
   U1403 : MUX2_X1 port map( A => n1103, B => n1041, S => n816, Z => n1009);
   U1404 : MUX2_X1 port map( A => n961, B => n1009, S => RF_RD2_DATA(4), Z => 
                           n962);
   U1405 : MUX2_X1 port map( A => n962, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN267);
   U1406 : MUX2_X1 port map( A => n964, B => n963, S => n820, Z => n1089);
   U1407 : MUX2_X1 port map( A => n966, B => n965, S => n820, Z => n997);
   U1408 : MUX2_X1 port map( A => n1089, B => n997, S => n818, Z => n1058);
   U1409 : MUX2_X1 port map( A => n968, B => n967, S => n820, Z => n996);
   U1410 : MUX2_X1 port map( A => n970, B => n969, S => n820, Z => n999);
   U1411 : MUX2_X1 port map( A => n996, B => n999, S => n818, Z => n1017);
   U1412 : MUX2_X1 port map( A => n1058, B => n1017, S => n816, Z => n974);
   U1413 : MUX2_X1 port map( A => n972, B => n971, S => n820, Z => n998);
   U1414 : MUX2_X1 port map( A => n973, B => n780, S => n820, Z => n1000);
   U1415 : MUX2_X1 port map( A => n998, B => n1000, S => n819, Z => n1016);
   U1416 : MUX2_X1 port map( A => n1016, B => n781, S => n816, Z => n1045);
   U1417 : MUX2_X1 port map( A => n974, B => n1045, S => RF_RD2_DATA(4), Z => 
                           n975);
   U1418 : MUX2_X1 port map( A => n975, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN277);
   U1419 : MUX2_X1 port map( A => RF_RD1_DATA(11), B => RF_RD1_DATA(12), S => 
                           n822, Z => n1024);
   U1420 : MUX2_X1 port map( A => RF_RD1_DATA(13), B => RF_RD1_DATA(14), S => 
                           n822, Z => n986);
   U1421 : MUX2_X1 port map( A => n1024, B => n986, S => n820, Z => n1096);
   U1422 : MUX2_X1 port map( A => RF_RD1_DATA(15), B => RF_RD1_DATA(16), S => 
                           n822, Z => n985);
   U1423 : MUX2_X1 port map( A => RF_RD1_DATA(17), B => RF_RD1_DATA(18), S => 
                           n823, Z => n988);
   U1424 : MUX2_X1 port map( A => n985, B => n988, S => n820, Z => n1004);
   U1425 : MUX2_X1 port map( A => n1096, B => n1004, S => n818, Z => n1070);
   U1426 : MUX2_X1 port map( A => RF_RD1_DATA(19), B => RF_RD1_DATA(20), S => 
                           n823, Z => n987);
   U1427 : MUX2_X1 port map( A => RF_RD1_DATA(21), B => RF_RD1_DATA(22), S => 
                           n823, Z => n990);
   U1428 : MUX2_X1 port map( A => n987, B => n990, S => n820, Z => n1003);
   U1429 : MUX2_X1 port map( A => RF_RD1_DATA(23), B => RF_RD1_DATA(24), S => 
                           n823, Z => n989);
   U1430 : MUX2_X1 port map( A => RF_RD1_DATA(25), B => RF_RD1_DATA(26), S => 
                           n823, Z => n992);
   U1431 : MUX2_X1 port map( A => n989, B => n992, S => n820, Z => n1006);
   U1432 : MUX2_X1 port map( A => n1003, B => n1006, S => n818, Z => n1020);
   U1433 : MUX2_X1 port map( A => n1070, B => n1020, S => n816, Z => n976);
   U1434 : MUX2_X1 port map( A => RF_RD1_DATA(27), B => RF_RD1_DATA(28), S => 
                           n823, Z => n991);
   U1435 : MUX2_X1 port map( A => RF_RD1_DATA(29), B => RF_RD1_DATA(30), S => 
                           n823, Z => n993);
   U1436 : MUX2_X1 port map( A => n991, B => n993, S => n820, Z => n1005);
   U1437 : MUX2_X1 port map( A => n1005, B => n780, S => n818, Z => n1019);
   U1438 : MUX2_X1 port map( A => n1019, B => n781, S => n816, Z => n1047);
   U1439 : MUX2_X1 port map( A => n976, B => n1047, S => RF_RD2_DATA(4), Z => 
                           n977);
   U1440 : MUX2_X1 port map( A => n977, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN278);
   U1441 : MUX2_X1 port map( A => n979, B => n978, S => n818, Z => n1077);
   U1442 : MUX2_X1 port map( A => n981, B => n980, S => n818, Z => n1031);
   U1443 : MUX2_X1 port map( A => n1077, B => n1031, S => n817, Z => n983);
   U1444 : MUX2_X1 port map( A => n982, B => n780, S => n818, Z => n1030);
   U1445 : MUX2_X1 port map( A => n1030, B => n781, S => n816, Z => n1049);
   U1446 : MUX2_X1 port map( A => n983, B => n1049, S => RF_RD2_DATA(4), Z => 
                           n984);
   U1447 : MUX2_X1 port map( A => n984, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN279);
   U1448 : MUX2_X1 port map( A => n986, B => n985, S => n821, Z => n1025);
   U1449 : MUX2_X1 port map( A => n988, B => n987, S => n821, Z => n1012);
   U1450 : MUX2_X1 port map( A => n1025, B => n1012, S => n818, Z => n1084);
   U1451 : MUX2_X1 port map( A => n990, B => n989, S => n821, Z => n1011);
   U1452 : MUX2_X1 port map( A => n992, B => n991, S => n821, Z => n1014);
   U1453 : MUX2_X1 port map( A => n1011, B => n1014, S => n818, Z => n1034);
   U1454 : MUX2_X1 port map( A => n1084, B => n1034, S => n816, Z => n994);
   U1455 : MUX2_X1 port map( A => n993, B => n780, S => n821, Z => n1013);
   U1456 : MUX2_X1 port map( A => n1013, B => n780, S => n819, Z => n1033);
   U1457 : MUX2_X1 port map( A => n1033, B => n781, S => n816, Z => n1051);
   U1458 : MUX2_X1 port map( A => n994, B => n1051, S => RF_RD2_DATA(4), Z => 
                           n995);
   U1459 : MUX2_X1 port map( A => n995, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN280);
   U1460 : MUX2_X1 port map( A => n997, B => n996, S => n819, Z => n1091);
   U1461 : MUX2_X1 port map( A => n999, B => n998, S => n819, Z => n1037);
   U1462 : MUX2_X1 port map( A => n1091, B => n1037, S => n816, Z => n1001);
   U1463 : MUX2_X1 port map( A => n1000, B => n781, S => n819, Z => n1036);
   U1464 : MUX2_X1 port map( A => n1036, B => n780, S => n816, Z => n1063);
   U1465 : MUX2_X1 port map( A => n1001, B => n1063, S => RF_RD2_DATA(4), Z => 
                           n1002);
   U1466 : MUX2_X1 port map( A => n1002, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(5), Z => DATAPATH_IxThird_stxALU1xN281);
   U1467 : MUX2_X1 port map( A => n1004, B => n1003, S => n819, Z => n1098);
   U1468 : MUX2_X1 port map( A => n1006, B => n1005, S => n819, Z => n1039);
   U1469 : MUX2_X1 port map( A => n1098, B => n1039, S => n816, Z => n1007);
   U1470 : MUX2_X1 port map( A => n1007, B => RF_RD1_DATA(31), S => 
                           RF_RD2_DATA(4), Z => n1008);
   U1471 : MUX2_X1 port map( A => n1008, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN282);
   U1472 : MUX2_X1 port map( A => n1009, B => n781, S => RF_RD2_DATA(4), Z => 
                           n1010);
   U1473 : MUX2_X1 port map( A => n1010, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN283);
   U1474 : MUX2_X1 port map( A => n1012, B => n1011, S => n819, Z => n1108);
   U1475 : MUX2_X1 port map( A => n1014, B => n1013, S => n819, Z => n1043);
   U1476 : MUX2_X1 port map( A => n1108, B => n1043, S => n816, Z => n1027);
   U1477 : MUX2_X1 port map( A => n1027, B => n781, S => RF_RD2_DATA(4), Z => 
                           n1015);
   U1478 : MUX2_X1 port map( A => n1015, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN284);
   U1479 : MUX2_X1 port map( A => n1017, B => n1016, S => n816, Z => n1060);
   U1480 : MUX2_X1 port map( A => n1060, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1018);
   U1481 : MUX2_X1 port map( A => n1018, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN285);
   U1482 : MUX2_X1 port map( A => n1020, B => n1019, S => n817, Z => n1072);
   U1483 : MUX2_X1 port map( A => n1072, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1021);
   U1484 : MUX2_X1 port map( A => n1021, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN286);
   U1485 : MUX2_X1 port map( A => RF_RD1_DATA(1), B => RF_RD1_DATA(2), S => 
                           n823, Z => n1022);
   U1486 : MUX2_X1 port map( A => RF_RD1_DATA(3), B => RF_RD1_DATA(4), S => 
                           n823, Z => n1066);
   U1487 : MUX2_X1 port map( A => n1022, B => n1066, S => n821, Z => n1023);
   U1488 : MUX2_X1 port map( A => RF_RD1_DATA(5), B => RF_RD1_DATA(6), S => 
                           n823, Z => n1065);
   U1489 : MUX2_X1 port map( A => RF_RD1_DATA(7), B => RF_RD1_DATA(8), S => 
                           n823, Z => n1068);
   U1490 : MUX2_X1 port map( A => n1065, B => n1068, S => n821, Z => n1083);
   U1491 : MUX2_X1 port map( A => n1023, B => n1083, S => n819, Z => n1026);
   U1492 : MUX2_X1 port map( A => RF_RD1_DATA(9), B => RF_RD1_DATA(10), S => 
                           n823, Z => n1067);
   U1493 : MUX2_X1 port map( A => n1067, B => n1024, S => n821, Z => n1082);
   U1494 : MUX2_X1 port map( A => n1082, B => n1025, S => n819, Z => n1109);
   U1495 : MUX2_X1 port map( A => n1026, B => n1109, S => n817, Z => n1028);
   U1496 : MUX2_X1 port map( A => n1028, B => n1027, S => RF_RD2_DATA(4), Z => 
                           n1029);
   U1497 : MUX2_X1 port map( A => n1029, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN268);
   U1498 : MUX2_X1 port map( A => n1031, B => n1030, S => n817, Z => n1079);
   U1499 : MUX2_X1 port map( A => n1079, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1032);
   U1500 : MUX2_X1 port map( A => n1032, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN287);
   U1501 : MUX2_X1 port map( A => n1034, B => n1033, S => n817, Z => n1086);
   U1502 : MUX2_X1 port map( A => n1086, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1035);
   U1503 : MUX2_X1 port map( A => n1035, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN288);
   U1504 : MUX2_X1 port map( A => n1037, B => n1036, S => n817, Z => n1093);
   U1505 : MUX2_X1 port map( A => n1093, B => n779, S => RF_RD2_DATA(4), Z => 
                           n1038);
   U1506 : MUX2_X1 port map( A => n1038, B => n779, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN289);
   U1507 : MUX2_X1 port map( A => n1039, B => n779, S => n817, Z => n1100);
   U1508 : MUX2_X1 port map( A => n1100, B => n779, S => RF_RD2_DATA(4), Z => 
                           n1040);
   U1509 : MUX2_X1 port map( A => n1040, B => n779, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN290);
   U1510 : MUX2_X1 port map( A => n1041, B => n779, S => n817, Z => n1105);
   U1511 : MUX2_X1 port map( A => n1105, B => n779, S => RF_RD2_DATA(4), Z => 
                           n1042);
   U1512 : MUX2_X1 port map( A => n1042, B => n779, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN291);
   U1513 : MUX2_X1 port map( A => n1043, B => n779, S => n817, Z => n1110);
   U1514 : MUX2_X1 port map( A => n1110, B => n779, S => RF_RD2_DATA(4), Z => 
                           n1044);
   U1515 : MUX2_X1 port map( A => n1044, B => n779, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN292);
   U1516 : MUX2_X1 port map( A => n1045, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1046);
   U1517 : MUX2_X1 port map( A => n1046, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN293);
   U1518 : MUX2_X1 port map( A => n1047, B => n781, S => RF_RD2_DATA(4), Z => 
                           n1048);
   U1519 : MUX2_X1 port map( A => n1048, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN294);
   U1520 : MUX2_X1 port map( A => n1049, B => n781, S => RF_RD2_DATA(4), Z => 
                           n1050);
   U1521 : MUX2_X1 port map( A => n1050, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN295);
   U1522 : MUX2_X1 port map( A => n1051, B => n781, S => RF_RD2_DATA(4), Z => 
                           n1052);
   U1523 : MUX2_X1 port map( A => n1052, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN296);
   U1524 : MUX2_X1 port map( A => n1054, B => n1053, S => n821, Z => n1057);
   U1525 : MUX2_X1 port map( A => n1056, B => n1055, S => n821, Z => n1090);
   U1526 : MUX2_X1 port map( A => n1057, B => n1090, S => n819, Z => n1059);
   U1527 : MUX2_X1 port map( A => n1059, B => n1058, S => n817, Z => n1061);
   U1528 : MUX2_X1 port map( A => n1061, B => n1060, S => RF_RD2_DATA(4), Z => 
                           n1062);
   U1529 : MUX2_X1 port map( A => n1062, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN269);
   U1530 : MUX2_X1 port map( A => n1063, B => n780, S => RF_RD2_DATA(4), Z => 
                           n1064);
   U1531 : MUX2_X1 port map( A => n1064, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN297);
   U1532 : MUX2_X1 port map( A => n1066, B => n1065, S => n821, Z => n1069);
   U1533 : MUX2_X1 port map( A => n1068, B => n1067, S => n821, Z => n1097);
   U1534 : MUX2_X1 port map( A => n1069, B => n1097, S => n819, Z => n1071);
   U1535 : MUX2_X1 port map( A => n1071, B => n1070, S => n817, Z => n1073);
   U1536 : MUX2_X1 port map( A => n1073, B => n1072, S => RF_RD2_DATA(4), Z => 
                           n1074);
   U1537 : MUX2_X1 port map( A => n1074, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN270);
   U1538 : MUX2_X1 port map( A => n1076, B => n1075, S => n819, Z => n1078);
   U1539 : MUX2_X1 port map( A => n1078, B => n1077, S => n817, Z => n1080);
   U1540 : MUX2_X1 port map( A => n1080, B => n1079, S => RF_RD2_DATA(4), Z => 
                           n1081);
   U1541 : MUX2_X1 port map( A => n1081, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN271);
   U1542 : MUX2_X1 port map( A => n1083, B => n1082, S => n819, Z => n1085);
   U1543 : MUX2_X1 port map( A => n1085, B => n1084, S => n817, Z => n1087);
   U1544 : MUX2_X1 port map( A => n1087, B => n1086, S => RF_RD2_DATA(4), Z => 
                           n1088);
   U1545 : MUX2_X1 port map( A => n1088, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN272);
   U1546 : MUX2_X1 port map( A => n1090, B => n1089, S => n819, Z => n1092);
   U1547 : MUX2_X1 port map( A => n1092, B => n1091, S => n817, Z => n1094);
   U1548 : MUX2_X1 port map( A => n1094, B => n1093, S => RF_RD2_DATA(4), Z => 
                           n1095);
   U1549 : MUX2_X1 port map( A => n1095, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN273);
   U1550 : MUX2_X1 port map( A => n1097, B => n1096, S => n819, Z => n1099);
   U1551 : MUX2_X1 port map( A => n1099, B => n1098, S => n817, Z => n1101);
   U1552 : MUX2_X1 port map( A => n1101, B => n1100, S => RF_RD2_DATA(4), Z => 
                           n1102);
   U1553 : MUX2_X1 port map( A => n1102, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN274);
   U1554 : MUX2_X1 port map( A => n1104, B => n1103, S => n817, Z => n1106);
   U1555 : MUX2_X1 port map( A => n1106, B => n1105, S => RF_RD2_DATA(4), Z => 
                           n1107);
   U1556 : MUX2_X1 port map( A => n1107, B => n781, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN275);
   U1557 : MUX2_X1 port map( A => n1109, B => n1108, S => n817, Z => n1111);
   U1558 : MUX2_X1 port map( A => n1111, B => n1110, S => RF_RD2_DATA(4), Z => 
                           n1112);
   U1559 : MUX2_X1 port map( A => n1112, B => n780, S => RF_RD2_DATA(5), Z => 
                           DATAPATH_IxThird_stxALU1xN276);

end SYN_RV32I_rtl;
